magic
tech scmos
timestamp 1741142099
<< nwell >>
rect -4 30 36 91
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
rect 23 8 25 12
<< ptransistor >>
rect 7 36 9 48
rect 12 36 14 48
rect 23 36 25 48
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
rect 14 8 15 12
rect 17 8 18 12
rect 22 8 23 12
rect 25 8 26 12
<< pdiffusion >>
rect 6 36 7 48
rect 9 36 12 48
rect 14 36 23 48
rect 25 36 26 48
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
rect 18 8 22 12
rect 26 8 30 12
<< pdcontact >>
rect 2 36 6 48
rect 26 36 30 48
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 84 6 88
<< polysilicon >>
rect 7 48 9 50
rect 12 48 14 50
rect 23 48 25 50
rect 7 12 9 36
rect 12 26 14 36
rect 23 33 25 36
rect 22 29 25 33
rect 16 22 17 26
rect 15 12 17 22
rect 23 12 25 29
rect 7 6 9 8
rect 15 6 17 8
rect 23 6 25 8
<< polycontact >>
rect 3 15 7 19
rect 18 29 22 33
rect 12 22 16 26
<< metal1 >>
rect 0 84 2 88
rect 6 84 32 88
rect 2 48 6 84
rect 0 29 18 33
rect 0 22 12 26
rect 26 19 30 36
rect 0 15 3 19
rect 10 15 30 19
rect 10 12 14 15
rect 26 12 30 15
rect 2 4 6 8
rect 18 4 22 8
rect 0 0 2 4
rect 6 0 32 4
<< labels >>
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel metal1 28 18 28 18 1 Y
rlabel metal1 2 17 2 17 1 A
rlabel metal1 2 24 2 24 1 B
rlabel metal1 2 31 2 31 1 C
rlabel nsubstratencontact 4 86 4 86 1 VDD
<< end >>
