magic
tech scmos
timestamp 1741221395
<< nwell >>
rect -5 70 38 91
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
rect 24 8 26 12
<< ptransistor >>
rect 7 76 9 80
rect 15 76 17 80
rect 24 76 26 80
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 15 12
rect 17 8 24 12
rect 26 8 27 12
<< pdiffusion >>
rect 6 76 7 80
rect 9 76 10 80
rect 14 76 15 80
rect 17 76 18 80
rect 22 76 24 80
rect 26 76 27 80
<< ndcontact >>
rect 2 8 6 12
rect 27 8 31 12
<< pdcontact >>
rect 2 76 6 80
rect 10 76 14 80
rect 18 76 22 80
rect 27 76 31 80
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 10 84 14 88
rect 27 84 31 88
<< polysilicon >>
rect 7 80 9 82
rect 15 80 17 82
rect 24 80 26 82
rect 7 12 9 76
rect 15 45 17 76
rect 16 41 17 45
rect 15 12 17 41
rect 24 12 26 76
rect 7 6 9 8
rect 15 6 17 8
rect 24 6 26 8
<< polycontact >>
rect 3 24 7 28
rect 20 58 24 62
rect 12 41 16 45
<< metal1 >>
rect 0 84 10 88
rect 14 84 27 88
rect 31 84 33 88
rect 10 80 14 84
rect 27 80 31 84
rect 2 72 6 76
rect 18 72 22 76
rect 2 68 31 72
rect 27 12 31 68
rect 2 4 6 8
rect 0 0 2 4
rect 6 0 33 4
<< labels >>
rlabel nsubstratencontact 12 86 12 86 1 VDD
rlabel nsubstratencontact 29 86 29 86 1 VDD
rlabel polycontact 5 26 5 26 1 A
rlabel polycontact 14 43 14 43 1 B
rlabel polycontact 22 60 22 60 1 C
rlabel metal1 29 34 29 34 1 Y
rlabel psubstratepcontact 4 2 4 2 1 VSS
<< end >>
