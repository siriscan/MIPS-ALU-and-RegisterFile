magic
tech scmos
timestamp 1746770961
<< metal1 >>
rect -803 332 -574 336
rect -63 332 16 336
rect -795 248 -574 252
rect -62 248 15 252
rect -785 240 -572 244
rect -785 224 14 228
rect -184 216 23 220
rect -785 200 -524 204
rect -512 200 -60 204
rect -56 200 0 204
rect 2930 200 2934 204
rect 2938 200 2994 204
rect -785 192 -460 196
rect -448 192 -52 196
rect -48 192 0 196
rect 2930 192 2942 196
rect 2946 192 2994 196
rect -785 184 -396 188
rect -384 184 -44 188
rect -40 184 0 188
rect 2930 184 2950 188
rect 2954 184 2994 188
rect -785 176 -332 180
rect -320 176 -36 180
rect -32 176 0 180
rect 2930 176 2958 180
rect 2962 176 2994 180
rect -785 168 -268 172
rect -256 168 -28 172
rect -24 168 0 172
rect 2930 168 2966 172
rect 2970 168 2994 172
rect -785 160 -204 164
rect -192 160 -20 164
rect -16 160 0 164
rect 2930 160 2974 164
rect 2978 160 2994 164
rect -785 152 -140 156
rect -128 152 -12 156
rect -8 152 0 156
rect 2930 152 2982 156
rect 2986 152 2994 156
rect -785 144 -76 148
rect -64 144 -4 148
rect 2930 144 2990 148
rect 2909 136 2925 140
rect 2909 128 2925 132
rect 2909 120 2925 124
rect 2909 112 2925 116
rect 2909 104 2925 108
rect 2909 96 2925 100
rect 2909 88 2925 92
rect 2909 80 2925 84
rect 2930 72 2998 76
rect 3002 72 3058 76
rect 2930 64 3006 68
rect 3010 64 3058 68
rect 2930 56 3014 60
rect 3018 56 3058 60
rect 2930 48 3022 52
rect 3026 48 3058 52
rect 2930 40 3030 44
rect 3034 40 3058 44
rect 2930 32 3038 36
rect 3042 32 3058 36
rect -74 24 6 28
rect 2930 24 3046 28
rect 3050 24 3058 28
rect -64 16 7 20
rect 2929 16 3054 20
rect -803 -8 -600 -4
rect -82 -8 14 -4
rect -795 -92 -600 -88
rect -82 -92 15 -88
rect -785 -100 -598 -96
rect -178 -100 14 -96
rect -785 -108 -578 -104
rect -785 -124 -566 -120
rect -785 -140 -550 -136
rect -56 -140 0 -136
rect 2930 -140 2934 -136
rect 2938 -140 2994 -136
rect -60 -148 -52 -144
rect -48 -148 0 -144
rect 2930 -148 2942 -144
rect 2946 -148 2994 -144
rect -60 -156 -44 -152
rect -40 -156 0 -152
rect 2930 -156 2950 -152
rect 2954 -156 2994 -152
rect -60 -164 -36 -160
rect -32 -164 0 -160
rect 2930 -164 2958 -160
rect 2962 -164 2994 -160
rect -60 -172 -28 -168
rect -24 -172 0 -168
rect 2930 -172 2966 -168
rect 2970 -172 2994 -168
rect -60 -180 -20 -176
rect -16 -180 0 -176
rect 2930 -180 2974 -176
rect 2978 -180 2994 -176
rect -60 -188 -12 -184
rect -8 -188 0 -184
rect 2930 -188 2982 -184
rect 2986 -188 2994 -184
rect -60 -196 -4 -192
rect 2930 -196 2990 -192
rect 2909 -204 2925 -200
rect 2909 -212 2925 -208
rect -465 -220 -78 -216
rect 2909 -220 2925 -216
rect -424 -228 -94 -224
rect 2909 -228 2925 -224
rect 2909 -236 2925 -232
rect -803 -243 -568 -239
rect -176 -243 -86 -239
rect 2909 -244 2925 -240
rect 2909 -252 2925 -248
rect 2909 -260 2925 -256
rect 2930 -268 2998 -264
rect 3002 -268 3058 -264
rect 2930 -276 3006 -272
rect 3010 -276 3058 -272
rect 2930 -284 3014 -280
rect 3018 -284 3058 -280
rect 2930 -292 3022 -288
rect 3026 -292 3058 -288
rect 2930 -300 3030 -296
rect 3034 -300 3058 -296
rect 2930 -308 3038 -304
rect 3042 -308 3058 -304
rect -90 -316 7 -312
rect 2930 -316 3046 -312
rect 3050 -316 3058 -312
rect -795 -327 -565 -323
rect -72 -324 6 -320
rect 2930 -324 3054 -320
rect -785 -343 -550 -339
rect -82 -348 14 -344
rect -785 -359 -534 -355
rect -785 -375 -518 -371
rect -371 -432 15 -428
rect -162 -440 36 -436
rect -684 -468 -68 -464
rect -643 -476 -76 -472
rect -56 -480 0 -476
rect 2930 -480 2934 -476
rect 2938 -480 2994 -476
rect -803 -491 -719 -487
rect -60 -488 -52 -484
rect -48 -488 0 -484
rect 2930 -488 2942 -484
rect 2946 -488 2994 -484
rect -60 -496 -44 -492
rect -40 -496 0 -492
rect 2930 -496 2950 -492
rect 2954 -496 2994 -492
rect -60 -504 -36 -500
rect -32 -504 0 -500
rect 2930 -504 2958 -500
rect 2962 -504 2994 -500
rect -60 -512 -28 -508
rect -24 -512 0 -508
rect 2930 -512 2966 -508
rect 2970 -512 2994 -508
rect -60 -520 -20 -516
rect -16 -520 0 -516
rect 2930 -520 2974 -516
rect 2978 -520 2994 -516
rect -60 -528 -12 -524
rect -8 -528 0 -524
rect 2930 -528 2982 -524
rect 2986 -528 2994 -524
rect -60 -536 -4 -532
rect 2930 -536 2990 -532
rect 2909 -544 2925 -540
rect 2909 -552 2925 -548
rect 2909 -560 2925 -556
rect 2909 -568 2925 -564
rect -795 -575 -786 -571
rect -396 -575 -375 -571
rect 2909 -576 2925 -572
rect 2909 -584 2925 -580
rect -785 -591 -769 -587
rect 2909 -592 2925 -588
rect 2909 -600 2925 -596
rect -785 -607 -753 -603
rect 2930 -608 2998 -604
rect 3002 -608 3058 -604
rect 2930 -616 3006 -612
rect 3010 -616 3058 -612
rect -785 -623 -737 -619
rect 2930 -624 3014 -620
rect 3018 -624 3058 -620
rect 2930 -632 3022 -628
rect 3026 -632 3058 -628
rect 2930 -640 3030 -636
rect 3034 -640 3058 -636
rect 2930 -648 3038 -644
rect 3042 -648 3058 -644
rect -383 -656 6 -652
rect 2930 -656 3046 -652
rect 3050 -656 3058 -652
rect -602 -664 6 -660
rect 2930 -664 3054 -660
rect -803 -688 14 -684
rect -795 -772 15 -768
rect -146 -780 14 -776
rect -56 -820 0 -816
rect 2930 -820 2934 -816
rect 2938 -820 2994 -816
rect -60 -828 -52 -824
rect -48 -828 0 -824
rect 2930 -828 2942 -824
rect 2946 -828 2994 -824
rect -60 -836 -44 -832
rect -40 -836 0 -832
rect 2930 -836 2950 -832
rect 2954 -836 2994 -832
rect -60 -844 -36 -840
rect -32 -844 0 -840
rect 2930 -844 2958 -840
rect 2962 -844 2994 -840
rect -60 -852 -28 -848
rect -24 -852 0 -848
rect 2930 -852 2966 -848
rect 2970 -852 2994 -848
rect -60 -860 -20 -856
rect -16 -860 0 -856
rect 2930 -860 2974 -856
rect 2978 -860 2994 -856
rect -60 -868 -12 -864
rect -8 -868 0 -864
rect 2930 -868 2982 -864
rect 2986 -868 2994 -864
rect -60 -876 -4 -872
rect 2930 -876 2990 -872
rect 2910 -884 2926 -880
rect 2910 -892 2926 -888
rect 2910 -900 2926 -896
rect 2910 -908 2926 -904
rect 2910 -916 2926 -912
rect 2910 -924 2926 -920
rect 2910 -932 2926 -928
rect 2910 -940 2926 -936
rect 2930 -948 2998 -944
rect 3002 -948 3058 -944
rect 2930 -956 3006 -952
rect 3010 -956 3058 -952
rect 2930 -964 3014 -960
rect 3018 -964 3058 -960
rect 2930 -972 3022 -968
rect 3026 -972 3058 -968
rect 2930 -980 3030 -976
rect 3034 -980 3058 -976
rect 2930 -988 3038 -984
rect 3042 -988 3058 -984
rect -342 -996 6 -992
rect 2930 -996 3046 -992
rect 3050 -996 3058 -992
rect -561 -1004 15 -1000
rect 2930 -1004 3054 -1000
rect -803 -1028 14 -1024
rect -795 -1112 15 -1108
rect -130 -1120 14 -1116
rect -56 -1160 0 -1156
rect 2930 -1160 2934 -1156
rect -60 -1168 -52 -1164
rect -48 -1168 0 -1164
rect 2930 -1168 2934 -1164
rect -60 -1176 -44 -1172
rect -40 -1176 0 -1172
rect 2930 -1176 2934 -1172
rect -60 -1184 -36 -1180
rect -32 -1184 0 -1180
rect 2930 -1184 2934 -1180
rect -60 -1192 -28 -1188
rect -24 -1192 0 -1188
rect 2930 -1192 2934 -1188
rect -60 -1200 -20 -1196
rect -16 -1200 0 -1196
rect 2930 -1200 2934 -1196
rect -60 -1208 -12 -1204
rect -8 -1208 0 -1204
rect 2930 -1208 2934 -1204
rect -60 -1216 -4 -1212
rect 2930 -1216 2934 -1212
rect 2910 -1224 2926 -1220
rect 2910 -1232 2926 -1228
rect 2910 -1240 2926 -1236
rect 2910 -1248 2926 -1244
rect 2910 -1256 2926 -1252
rect 2910 -1264 2926 -1260
rect 2910 -1272 2926 -1268
rect 2910 -1280 2926 -1276
rect 2930 -1288 2998 -1284
rect 3002 -1288 3058 -1284
rect 2930 -1296 3006 -1292
rect 3010 -1296 3058 -1292
rect 2930 -1304 3014 -1300
rect 3018 -1304 3058 -1300
rect 2930 -1312 3022 -1308
rect 3026 -1312 3058 -1308
rect 2930 -1320 3030 -1316
rect 3034 -1320 3058 -1316
rect 2930 -1328 3038 -1324
rect 3042 -1328 3058 -1324
rect -301 -1336 6 -1332
rect 2930 -1336 3046 -1332
rect 3050 -1336 3058 -1332
rect -520 -1344 6 -1340
rect 2930 -1344 3054 -1340
rect -803 -1368 14 -1364
rect -795 -1452 15 -1448
rect -114 -1460 14 -1456
rect -56 -1500 0 -1496
rect 2930 -1500 2934 -1496
rect 2938 -1500 2994 -1496
rect -60 -1508 -52 -1504
rect -48 -1508 0 -1504
rect 2930 -1508 2942 -1504
rect 2946 -1508 2994 -1504
rect -60 -1516 -44 -1512
rect -40 -1516 0 -1512
rect 2930 -1516 2950 -1512
rect 2954 -1516 2994 -1512
rect -60 -1524 -36 -1520
rect -32 -1524 0 -1520
rect 2930 -1524 2958 -1520
rect 2962 -1524 2994 -1520
rect -60 -1532 -28 -1528
rect -24 -1532 0 -1528
rect 2930 -1532 2966 -1528
rect 2970 -1532 2994 -1528
rect -60 -1540 -20 -1536
rect -16 -1540 0 -1536
rect 2930 -1540 2974 -1536
rect 2978 -1540 2994 -1536
rect -60 -1548 -12 -1544
rect -8 -1548 0 -1544
rect 2930 -1548 2982 -1544
rect 2986 -1548 2994 -1544
rect -60 -1556 -4 -1552
rect 2930 -1556 2990 -1552
rect 2910 -1564 2926 -1560
rect 2910 -1572 2926 -1568
rect 2910 -1580 2926 -1576
rect 2910 -1588 2926 -1584
rect 2910 -1596 2926 -1592
rect 2910 -1604 2926 -1600
rect 2910 -1612 2926 -1608
rect 2910 -1620 2926 -1616
rect 2930 -1628 2998 -1624
rect 3002 -1628 3058 -1624
rect 2930 -1636 3006 -1632
rect 3010 -1636 3058 -1632
rect 2930 -1644 3014 -1640
rect 3018 -1644 3058 -1640
rect 2930 -1652 3022 -1648
rect 3026 -1652 3058 -1648
rect 2930 -1660 3030 -1656
rect 3034 -1660 3058 -1656
rect 2930 -1668 3038 -1664
rect 3042 -1668 3058 -1664
rect -260 -1676 6 -1672
rect 2930 -1676 3046 -1672
rect 3050 -1676 3058 -1672
rect -479 -1684 6 -1680
rect 2930 -1684 3054 -1680
rect -803 -1708 14 -1704
rect -795 -1792 15 -1788
rect -98 -1800 39 -1796
rect -56 -1840 0 -1836
rect 2930 -1840 2934 -1836
rect 2938 -1840 2994 -1836
rect -60 -1848 -52 -1844
rect -48 -1848 0 -1844
rect 2930 -1848 2942 -1844
rect 2946 -1848 2994 -1844
rect -60 -1856 -44 -1852
rect -40 -1856 0 -1852
rect 2930 -1856 2950 -1852
rect 2954 -1856 2994 -1852
rect -60 -1864 -36 -1860
rect -32 -1864 0 -1860
rect 2930 -1864 2958 -1860
rect 2962 -1864 2994 -1860
rect -60 -1872 -28 -1868
rect -24 -1872 0 -1868
rect 2930 -1872 2966 -1868
rect 2970 -1872 2994 -1868
rect -60 -1880 -20 -1876
rect -16 -1880 0 -1876
rect 2930 -1880 2974 -1876
rect 2978 -1880 2994 -1876
rect -60 -1888 -12 -1884
rect -8 -1888 0 -1884
rect 2930 -1888 2982 -1884
rect 2986 -1888 2994 -1884
rect -60 -1896 -4 -1892
rect 2930 -1896 2990 -1892
rect 2910 -1904 2926 -1900
rect 2910 -1912 2926 -1908
rect 2910 -1920 2926 -1916
rect 2910 -1928 2926 -1924
rect 2910 -1936 2926 -1932
rect 2910 -1944 2926 -1940
rect 2910 -1952 2926 -1948
rect 2910 -1960 2926 -1956
rect 2930 -1968 2998 -1964
rect 3002 -1968 3058 -1964
rect 2930 -1976 3006 -1972
rect 3010 -1976 3058 -1972
rect 2930 -1984 3014 -1980
rect 3018 -1984 3058 -1980
rect 2930 -1992 3022 -1988
rect 3026 -1992 3058 -1988
rect 2930 -2000 3030 -1996
rect 3034 -2000 3058 -1996
rect 2930 -2008 3038 -2004
rect 3042 -2008 3058 -2004
rect -219 -2016 6 -2012
rect 2930 -2016 3046 -2012
rect 3050 -2016 3058 -2012
rect -438 -2024 6 -2020
rect 2930 -2024 3054 -2020
rect -803 -2040 -158 -2036
rect -795 -2124 -156 -2120
rect -178 -2132 -155 -2128
rect -397 -2140 -149 -2136
rect 732 -2148 2934 -2144
rect 2938 -2148 2994 -2144
rect 732 -2156 2942 -2152
rect 2946 -2156 2994 -2152
rect 732 -2164 2950 -2160
rect 2954 -2164 2994 -2160
rect 732 -2172 2958 -2168
rect 2962 -2172 2994 -2168
rect 732 -2180 2966 -2176
rect 2970 -2180 2994 -2176
rect 732 -2188 2974 -2184
rect 2978 -2188 2994 -2184
rect 732 -2196 2982 -2192
rect 2986 -2196 2994 -2192
rect 732 -2204 2990 -2200
rect 732 -2212 2926 -2208
rect 732 -2220 2998 -2216
rect 3002 -2220 3058 -2216
rect 732 -2228 3006 -2224
rect 3010 -2228 3058 -2224
rect 732 -2236 3014 -2232
rect 3018 -2236 3058 -2232
rect 732 -2244 3022 -2240
rect 3026 -2244 3058 -2240
rect 732 -2252 3030 -2248
rect 3034 -2252 3058 -2248
rect 732 -2260 3038 -2256
rect 3042 -2260 3058 -2256
rect 732 -2268 3046 -2264
rect 3050 -2268 3058 -2264
rect 732 -2276 3054 -2272
<< m2contact >>
rect -807 332 -803 336
rect -549 311 -545 315
rect -485 311 -481 315
rect -421 311 -417 315
rect -357 311 -353 315
rect -293 311 -289 315
rect -229 311 -225 315
rect -165 311 -161 315
rect -101 311 -97 315
rect -799 248 -795 252
rect 15 224 19 228
rect -188 216 -184 220
rect 23 216 27 220
rect -524 200 -520 204
rect -516 200 -512 204
rect -60 200 -56 204
rect 2934 200 2938 204
rect -460 192 -456 196
rect -452 192 -448 196
rect -52 192 -48 196
rect 2942 192 2946 196
rect -396 184 -392 188
rect -388 184 -384 188
rect -44 184 -40 188
rect 2950 184 2954 188
rect -332 176 -328 180
rect -324 176 -320 180
rect -36 176 -32 180
rect 2958 176 2962 180
rect -268 168 -264 172
rect -260 168 -256 172
rect -28 168 -24 172
rect 2966 168 2970 172
rect -204 160 -200 164
rect -196 160 -192 164
rect -20 160 -16 164
rect 2974 160 2978 164
rect -140 152 -136 156
rect -132 152 -128 156
rect -12 152 -8 156
rect 2982 152 2986 156
rect -76 144 -72 148
rect -68 144 -64 148
rect -4 144 0 148
rect 2990 144 2994 148
rect 2998 72 3002 76
rect 3006 64 3010 68
rect 3014 56 3018 60
rect 3022 48 3026 52
rect 3030 40 3034 44
rect 3038 32 3042 36
rect -78 24 -74 28
rect 3046 24 3050 28
rect -68 16 -64 20
rect 3054 16 3058 20
rect -807 -8 -803 -4
rect -799 -92 -795 -88
rect -598 -100 -594 -96
rect -182 -100 -178 -96
rect 15 -116 19 -112
rect -60 -140 -56 -136
rect 2934 -140 2938 -136
rect -52 -148 -48 -144
rect 2942 -148 2946 -144
rect -44 -156 -40 -152
rect 2950 -156 2954 -152
rect -36 -164 -32 -160
rect 2958 -164 2962 -160
rect -28 -172 -24 -168
rect 2966 -172 2970 -168
rect -20 -180 -16 -176
rect 2974 -180 2978 -176
rect -12 -188 -8 -184
rect 2982 -188 2986 -184
rect -4 -196 0 -192
rect 2990 -196 2994 -192
rect -469 -220 -465 -216
rect -78 -220 -74 -216
rect -428 -228 -424 -224
rect -94 -228 -90 -224
rect -807 -243 -803 -239
rect -86 -243 -82 -239
rect 2998 -268 3002 -264
rect 3006 -276 3010 -272
rect 3014 -284 3018 -280
rect 3022 -292 3026 -288
rect 3030 -300 3034 -296
rect 3038 -308 3042 -304
rect -94 -316 -90 -312
rect 3046 -316 3050 -312
rect -799 -327 -795 -323
rect -76 -324 -72 -320
rect 3054 -324 3058 -320
rect -566 -331 -562 -327
rect -86 -348 -82 -344
rect -375 -432 -371 -428
rect -166 -440 -162 -436
rect 15 -456 19 -452
rect -688 -468 -684 -464
rect -68 -468 -64 -464
rect -647 -476 -643 -472
rect -76 -476 -72 -472
rect -60 -480 -56 -476
rect 2934 -480 2938 -476
rect -807 -491 -803 -487
rect -52 -488 -48 -484
rect 2942 -488 2946 -484
rect -44 -496 -40 -492
rect 2950 -496 2954 -492
rect -36 -504 -32 -500
rect 2958 -504 2962 -500
rect -28 -512 -24 -508
rect 2966 -512 2970 -508
rect -20 -520 -16 -516
rect 2974 -520 2978 -516
rect -12 -528 -8 -524
rect 2982 -528 2986 -524
rect -4 -536 0 -532
rect 2990 -536 2994 -532
rect -799 -575 -795 -571
rect -375 -575 -371 -571
rect -785 -579 -781 -575
rect 2998 -608 3002 -604
rect 3006 -616 3010 -612
rect 3014 -624 3018 -620
rect 3022 -632 3026 -628
rect 3030 -640 3034 -636
rect 3038 -648 3042 -644
rect -387 -656 -383 -652
rect 3046 -656 3050 -652
rect -606 -664 -602 -660
rect 3054 -664 3058 -660
rect -807 -688 -803 -684
rect -799 -772 -795 -768
rect -150 -780 -146 -776
rect 15 -796 19 -792
rect -60 -820 -56 -816
rect 2934 -820 2938 -816
rect -52 -828 -48 -824
rect 2942 -828 2946 -824
rect -44 -836 -40 -832
rect 2950 -836 2954 -832
rect -36 -844 -32 -840
rect 2958 -844 2962 -840
rect -28 -852 -24 -848
rect 2966 -852 2970 -848
rect -20 -860 -16 -856
rect 2974 -860 2978 -856
rect -12 -868 -8 -864
rect 2982 -868 2986 -864
rect -4 -876 0 -872
rect 2990 -876 2994 -872
rect 2998 -948 3002 -944
rect 3006 -956 3010 -952
rect 3014 -964 3018 -960
rect 3022 -972 3026 -968
rect 3030 -980 3034 -976
rect 3038 -988 3042 -984
rect -346 -996 -342 -992
rect 3046 -996 3050 -992
rect -565 -1004 -561 -1000
rect 3054 -1004 3058 -1000
rect -807 -1028 -803 -1024
rect -799 -1112 -795 -1108
rect -134 -1120 -130 -1116
rect 15 -1136 19 -1132
rect -60 -1160 -56 -1156
rect -52 -1168 -48 -1164
rect -44 -1176 -40 -1172
rect -36 -1184 -32 -1180
rect -28 -1192 -24 -1188
rect -20 -1200 -16 -1196
rect -12 -1208 -8 -1204
rect -4 -1216 0 -1212
rect 2998 -1288 3002 -1284
rect 3006 -1296 3010 -1292
rect 3014 -1304 3018 -1300
rect 3022 -1312 3026 -1308
rect 3030 -1320 3034 -1316
rect 3038 -1328 3042 -1324
rect -305 -1336 -301 -1332
rect 3046 -1336 3050 -1332
rect -524 -1344 -520 -1340
rect 3054 -1344 3058 -1340
rect -807 -1368 -803 -1364
rect -799 -1452 -795 -1448
rect -118 -1460 -114 -1456
rect 15 -1476 19 -1472
rect -60 -1500 -56 -1496
rect 2934 -1500 2938 -1496
rect -52 -1508 -48 -1504
rect 2942 -1508 2946 -1504
rect -44 -1516 -40 -1512
rect 2950 -1516 2954 -1512
rect -36 -1524 -32 -1520
rect 2958 -1524 2962 -1520
rect -28 -1532 -24 -1528
rect 2966 -1532 2970 -1528
rect -20 -1540 -16 -1536
rect 2974 -1540 2978 -1536
rect -12 -1548 -8 -1544
rect 2982 -1548 2986 -1544
rect -4 -1556 0 -1552
rect 2990 -1556 2994 -1552
rect 2998 -1628 3002 -1624
rect 3006 -1636 3010 -1632
rect 3014 -1644 3018 -1640
rect 3022 -1652 3026 -1648
rect 3030 -1660 3034 -1656
rect 3038 -1668 3042 -1664
rect -264 -1676 -260 -1672
rect 3046 -1676 3050 -1672
rect -483 -1684 -479 -1680
rect 3054 -1684 3058 -1680
rect -807 -1708 -803 -1704
rect -799 -1792 -795 -1788
rect -102 -1800 -98 -1796
rect 15 -1816 19 -1812
rect -60 -1840 -56 -1836
rect 2934 -1840 2938 -1836
rect -52 -1848 -48 -1844
rect 2942 -1848 2946 -1844
rect -44 -1856 -40 -1852
rect 2950 -1856 2954 -1852
rect -36 -1864 -32 -1860
rect 2958 -1864 2962 -1860
rect -28 -1872 -24 -1868
rect 2966 -1872 2970 -1868
rect -20 -1880 -16 -1876
rect 2974 -1880 2978 -1876
rect -12 -1888 -8 -1884
rect 2982 -1888 2986 -1884
rect -4 -1896 0 -1892
rect 2990 -1896 2994 -1892
rect 2998 -1968 3002 -1964
rect 3006 -1976 3010 -1972
rect 3014 -1984 3018 -1980
rect 3022 -1992 3026 -1988
rect 3030 -2000 3034 -1996
rect 3038 -2008 3042 -2004
rect -223 -2016 -219 -2012
rect 3046 -2016 3050 -2012
rect -442 -2024 -438 -2020
rect 3054 -2024 3058 -2020
rect -807 -2040 -803 -2036
rect -799 -2124 -795 -2120
rect 86 -2124 90 -2120
rect -182 -2132 -178 -2128
rect -401 -2140 -397 -2136
rect 2934 -2148 2938 -2144
rect 2942 -2156 2946 -2152
rect 2950 -2164 2954 -2160
rect 2958 -2172 2962 -2168
rect 2966 -2180 2970 -2176
rect 2974 -2188 2978 -2184
rect 2982 -2196 2986 -2192
rect 2990 -2204 2994 -2200
rect 2998 -2220 3002 -2216
rect 3006 -2228 3010 -2224
rect 3014 -2236 3018 -2232
rect 3022 -2244 3026 -2240
rect 3030 -2252 3034 -2248
rect 3038 -2260 3042 -2256
rect 3046 -2268 3050 -2264
rect 3054 -2276 3058 -2272
<< metal2 >>
rect -807 -4 -803 332
rect -549 315 -545 345
rect -485 315 -481 345
rect -421 315 -417 345
rect -357 315 -353 345
rect -293 315 -289 345
rect -229 315 -225 345
rect -165 315 -161 345
rect -101 315 -97 345
rect -807 -239 -803 -8
rect -807 -487 -803 -243
rect -807 -684 -803 -491
rect -807 -1024 -803 -688
rect -807 -1364 -803 -1028
rect -807 -1704 -803 -1368
rect -807 -2036 -803 -1708
rect -799 -88 -795 248
rect -524 204 -520 288
rect -516 204 -512 232
rect -460 196 -456 288
rect -452 196 -448 232
rect -396 188 -392 288
rect -388 188 -384 232
rect -332 180 -328 288
rect -324 180 -320 232
rect -268 172 -264 288
rect -260 172 -256 232
rect -204 164 -200 288
rect -196 164 -192 232
rect -188 7 -184 216
rect -140 156 -136 288
rect -132 156 -128 232
rect -76 148 -72 288
rect -68 148 -64 232
rect -198 3 -184 7
rect -198 -76 -194 3
rect -799 -323 -795 -92
rect -469 -312 -465 -220
rect -428 -311 -424 -228
rect -799 -571 -795 -327
rect -688 -563 -684 -468
rect -647 -563 -643 -476
rect -799 -768 -795 -575
rect -606 -660 -602 -638
rect -799 -1108 -795 -772
rect -565 -1000 -561 -639
rect -799 -1448 -795 -1112
rect -524 -1340 -520 -639
rect -799 -1788 -795 -1452
rect -483 -1680 -479 -639
rect -799 -2120 -795 -1792
rect -442 -2020 -438 -639
rect -401 -2136 -397 -639
rect -387 -652 -383 -391
rect -375 -571 -371 -432
rect -346 -992 -342 -391
rect -305 -1332 -301 -391
rect -264 -1672 -260 -391
rect -223 -2012 -219 -391
rect -182 -2128 -178 -391
rect -166 -436 -162 -80
rect -150 -776 -146 -100
rect -134 -1116 -130 -100
rect -118 -1456 -114 -100
rect -102 -1796 -98 -84
rect -86 -109 -82 -100
rect -78 -216 -74 24
rect -94 -312 -90 -228
rect -86 -344 -82 -243
rect -76 -472 -72 -324
rect -68 -464 -64 16
rect -60 -136 -56 200
rect -60 -476 -56 -140
rect -60 -816 -56 -480
rect -60 -1156 -56 -820
rect -60 -1496 -56 -1160
rect -60 -1836 -56 -1500
rect -60 -1896 -56 -1840
rect -52 -144 -48 192
rect -52 -484 -48 -148
rect -52 -824 -48 -488
rect -52 -1164 -48 -828
rect -52 -1504 -48 -1168
rect -52 -1844 -48 -1508
rect -52 -1896 -48 -1848
rect -44 -152 -40 184
rect -44 -492 -40 -156
rect -44 -832 -40 -496
rect -44 -1172 -40 -836
rect -44 -1512 -40 -1176
rect -44 -1852 -40 -1516
rect -44 -1896 -40 -1856
rect -36 -160 -32 176
rect -36 -500 -32 -164
rect -36 -840 -32 -504
rect -36 -1180 -32 -844
rect -36 -1520 -32 -1184
rect -36 -1860 -32 -1524
rect -36 -1896 -32 -1864
rect -28 -168 -24 168
rect -28 -508 -24 -172
rect -28 -848 -24 -512
rect -28 -1188 -24 -852
rect -28 -1528 -24 -1192
rect -28 -1868 -24 -1532
rect -28 -1896 -24 -1872
rect -20 -176 -16 160
rect -20 -516 -16 -180
rect -20 -856 -16 -520
rect -20 -1196 -16 -860
rect -20 -1536 -16 -1200
rect -20 -1876 -16 -1540
rect -20 -1896 -16 -1880
rect -12 -184 -8 152
rect -12 -524 -8 -188
rect -12 -864 -8 -528
rect -12 -1204 -8 -868
rect -12 -1544 -8 -1208
rect -12 -1884 -8 -1548
rect -12 -1896 -8 -1888
rect -4 -192 0 144
rect -4 -532 0 -196
rect -4 -872 0 -536
rect -4 -1212 0 -876
rect -4 -1552 0 -1216
rect -4 -1892 0 -1556
rect 15 -112 19 224
rect 23 220 27 240
rect 15 -452 19 -116
rect 15 -792 19 -456
rect 15 -1132 19 -796
rect 15 -1472 19 -1136
rect 15 -1812 19 -1476
rect 2934 204 2938 220
rect 2934 -136 2938 200
rect 2934 -476 2938 -140
rect 2934 -816 2938 -480
rect 2934 -1496 2938 -820
rect 2934 -1836 2938 -1500
rect 2934 -2144 2938 -1840
rect 2934 -2276 2938 -2148
rect 2942 196 2946 220
rect 2942 -144 2946 192
rect 2942 -484 2946 -148
rect 2942 -824 2946 -488
rect 2942 -1504 2946 -828
rect 2942 -1844 2946 -1508
rect 2942 -2152 2946 -1848
rect 2942 -2276 2946 -2156
rect 2950 188 2954 220
rect 2950 -152 2954 184
rect 2950 -492 2954 -156
rect 2950 -832 2954 -496
rect 2950 -1512 2954 -836
rect 2950 -1852 2954 -1516
rect 2950 -2160 2954 -1856
rect 2950 -2276 2954 -2164
rect 2958 180 2962 220
rect 2958 -160 2962 176
rect 2958 -500 2962 -164
rect 2958 -840 2962 -504
rect 2958 -1520 2962 -844
rect 2958 -1860 2962 -1524
rect 2958 -2168 2962 -1864
rect 2958 -2276 2962 -2172
rect 2966 172 2970 220
rect 2966 -168 2970 168
rect 2966 -508 2970 -172
rect 2966 -848 2970 -512
rect 2966 -1528 2970 -852
rect 2966 -1868 2970 -1532
rect 2966 -2176 2970 -1872
rect 2966 -2276 2970 -2180
rect 2974 164 2978 220
rect 2974 -176 2978 160
rect 2974 -516 2978 -180
rect 2974 -856 2978 -520
rect 2974 -1536 2978 -860
rect 2974 -1876 2978 -1540
rect 2974 -2184 2978 -1880
rect 2974 -2276 2978 -2188
rect 2982 156 2986 220
rect 2982 -184 2986 152
rect 2982 -524 2986 -188
rect 2982 -864 2986 -528
rect 2982 -1544 2986 -868
rect 2982 -1884 2986 -1548
rect 2982 -2192 2986 -1888
rect 2982 -2276 2986 -2196
rect 2990 148 2994 220
rect 2990 -192 2994 144
rect 2990 -532 2994 -196
rect 2990 -872 2994 -536
rect 2990 -1552 2994 -876
rect 2990 -1892 2994 -1556
rect 2990 -2200 2994 -1896
rect 2990 -2276 2994 -2204
rect 2998 76 3002 220
rect 2998 -264 3002 72
rect 2998 -604 3002 -268
rect 2998 -944 3002 -608
rect 2998 -1284 3002 -948
rect 2998 -1624 3002 -1288
rect 2998 -1964 3002 -1628
rect 2998 -2216 3002 -1968
rect 2998 -2276 3002 -2220
rect 3006 68 3010 220
rect 3006 -272 3010 64
rect 3006 -612 3010 -276
rect 3006 -952 3010 -616
rect 3006 -1292 3010 -956
rect 3006 -1632 3010 -1296
rect 3006 -1972 3010 -1636
rect 3006 -2224 3010 -1976
rect 3006 -2276 3010 -2228
rect 3014 60 3018 220
rect 3014 -280 3018 56
rect 3014 -620 3018 -284
rect 3014 -960 3018 -624
rect 3014 -1300 3018 -964
rect 3014 -1640 3018 -1304
rect 3014 -1980 3018 -1644
rect 3014 -2232 3018 -1984
rect 3014 -2276 3018 -2236
rect 3022 52 3026 220
rect 3022 -288 3026 48
rect 3022 -628 3026 -292
rect 3022 -968 3026 -632
rect 3022 -1308 3026 -972
rect 3022 -1648 3026 -1312
rect 3022 -1988 3026 -1652
rect 3022 -2240 3026 -1992
rect 3022 -2276 3026 -2244
rect 3030 44 3034 220
rect 3030 -296 3034 40
rect 3030 -636 3034 -300
rect 3030 -976 3034 -640
rect 3030 -1316 3034 -980
rect 3030 -1656 3034 -1320
rect 3030 -1996 3034 -1660
rect 3030 -2248 3034 -2000
rect 3030 -2276 3034 -2252
rect 3038 36 3042 220
rect 3038 -304 3042 32
rect 3038 -644 3042 -308
rect 3038 -984 3042 -648
rect 3038 -1324 3042 -988
rect 3038 -1664 3042 -1328
rect 3038 -2004 3042 -1668
rect 3038 -2256 3042 -2008
rect 3038 -2276 3042 -2260
rect 3046 28 3050 220
rect 3046 -312 3050 24
rect 3046 -652 3050 -316
rect 3046 -992 3050 -656
rect 3046 -1332 3050 -996
rect 3046 -1672 3050 -1336
rect 3046 -2012 3050 -1676
rect 3046 -2264 3050 -2016
rect 3046 -2276 3050 -2268
rect 3054 20 3058 220
rect 3054 -320 3058 16
rect 3054 -660 3058 -324
rect 3054 -1000 3058 -664
rect 3054 -1340 3058 -1004
rect 3054 -1680 3058 -1344
rect 3054 -2020 3058 -1684
rect 3054 -2272 3058 -2024
use 8bitMUX2to1  8bitMUX2to1_0
timestamp 1746042099
transform 1 0 -578 0 1 232
box 0 0 520 107
use Decoder_4x8  Decoder_4x8_0
timestamp 1742681920
transform 1 0 -508 0 1 -327
box -64 -64 336 95
use Decoder_4x8  Decoder_4x8_1
timestamp 1742681920
transform 1 0 -727 0 1 -575
box -64 -64 336 95
use Decoder_Inv_4x8  Decoder_Inv_4x8_0
timestamp 1743018986
transform 1 0 -604 0 1 -156
box 0 -56 528 159
use REG0v2  REG0v2_0
timestamp 1746602637
transform 1 0 -158 0 1 -2136
box 0 -140 894 108
use REG8v2  REG8v2_0
timestamp 1746597901
transform 1 0 6 0 1 80
box -6 -64 2924 264
use REG8v2  REG8v2_1
timestamp 1746597901
transform 1 0 6 0 1 -260
box -6 -64 2924 264
use REG8v2  REG8v2_2
timestamp 1746597901
transform 1 0 6 0 1 -600
box -6 -64 2924 264
use REG8v2  REG8v2_3
timestamp 1746597901
transform 1 0 6 0 1 -940
box -6 -64 2924 264
use REG8v2  REG8v2_4
timestamp 1746597901
transform 1 0 6 0 1 -1280
box -6 -64 2924 264
use REG8v2  REG8v2_5
timestamp 1746597901
transform 1 0 6 0 1 -1620
box -6 -64 2924 264
use REG8v2  REG8v2_6
timestamp 1746597901
transform 1 0 6 0 1 -1960
box -6 -64 2924 264
<< labels >>
rlabel metal1 2922 138 2922 138 1 reg_zero0
rlabel metal1 2922 130 2922 130 1 reg_zero1
rlabel metal1 2922 122 2922 122 1 reg_zero2
rlabel metal1 2922 114 2922 114 1 reg_zero3
rlabel metal1 2922 106 2922 106 1 reg_zero4
rlabel metal1 2922 98 2922 98 1 reg_zero5
rlabel metal1 2922 90 2922 90 1 reg_zero6
rlabel metal1 2922 82 2922 82 1 reg_zero7
rlabel metal1 2925 -202 2925 -202 1 reg_one0
rlabel metal1 2925 -210 2925 -210 1 reg_one1
rlabel metal1 2925 -218 2925 -218 1 reg_one2
rlabel metal1 2925 -226 2925 -226 1 reg_one3
rlabel metal1 2925 -234 2925 -234 1 reg_one4
rlabel metal1 2925 -242 2925 -242 1 reg_one5
rlabel metal1 2925 -250 2925 -250 1 reg_one6
rlabel metal1 2925 -258 2925 -258 1 reg_one7
rlabel metal1 2925 -542 2925 -542 1 reg_two0
rlabel metal1 2925 -550 2925 -550 1 reg_two1
rlabel metal1 2925 -558 2925 -558 1 reg_two2
rlabel metal1 2925 -566 2925 -566 1 reg_two3
rlabel metal1 2924 -574 2924 -574 1 reg_two4
rlabel metal1 2925 -582 2925 -582 1 reg_two5
rlabel metal1 2925 -590 2925 -590 1 reg_two6
rlabel metal1 2925 -598 2925 -598 1 reg_two7
rlabel metal1 2924 -882 2924 -882 1 reg_three0
rlabel metal1 2924 -890 2924 -890 1 reg_three1
rlabel metal1 2924 -898 2924 -898 1 reg_three2
rlabel metal1 2924 -906 2924 -906 1 reg_three3
rlabel metal1 2924 -914 2924 -914 1 reg_three4
rlabel metal1 2924 -922 2924 -922 1 reg_three5
rlabel metal1 2924 -930 2924 -930 1 reg_three6
rlabel metal1 2924 -938 2924 -938 1 reg_three7
rlabel metal1 2925 -1222 2925 -1222 1 reg_four0
rlabel metal1 2925 -1230 2925 -1230 1 reg_four1
rlabel metal1 2925 -1238 2925 -1238 1 reg_four2
rlabel metal1 2925 -1246 2925 -1246 1 reg_four3
rlabel metal1 2925 -1254 2925 -1254 1 reg_four4
rlabel metal1 2925 -1262 2925 -1262 1 reg_four5
rlabel metal1 2926 -1270 2926 -1270 1 reg_four6
rlabel metal1 2926 -1278 2926 -1278 1 reg_four7
rlabel metal1 2926 -1562 2926 -1562 1 reg_five0
rlabel metal1 2926 -1570 2926 -1570 1 reg_five1
rlabel metal1 2925 -1578 2925 -1578 1 reg_five2
rlabel metal1 2925 -1586 2925 -1586 1 reg_five3
rlabel metal1 2925 -1594 2925 -1594 1 reg_five4
rlabel metal1 2925 -1602 2925 -1602 1 reg_five5
rlabel metal1 2925 -1610 2925 -1610 1 reg_five6
rlabel metal1 2925 -1618 2925 -1618 1 reg_five7
rlabel metal1 2923 -1902 2923 -1902 1 reg_six0
rlabel metal1 2923 -1910 2923 -1910 1 reg_six1
rlabel metal1 2923 -1918 2923 -1918 1 reg_six2
rlabel metal1 2923 -1926 2923 -1926 1 reg_six3
rlabel metal1 2923 -1934 2923 -1934 1 reg_six4
rlabel metal1 2923 -1942 2923 -1942 1 reg_six5
rlabel metal1 2923 -1950 2923 -1950 1 reg_six6
rlabel metal1 2923 -1958 2923 -1958 1 reg_six7
rlabel metal1 -782 -589 -782 -589 1 B_sel0
rlabel metal1 -782 -605 -782 -605 1 B_sel1
rlabel metal1 -782 -621 -782 -621 1 B_sel2
rlabel metal1 -782 -341 -782 -341 1 A_sel0
rlabel metal1 -782 -357 -782 -357 1 A_sel1
rlabel metal1 -782 -373 -782 -373 1 A_sel2
rlabel metal1 -781 -98 -781 -98 1 C_sel3
rlabel metal1 -781 -106 -781 -106 1 C_sel0
rlabel metal1 -781 -122 -781 -122 1 C_sel1
rlabel metal1 -782 -138 -782 -138 1 C_sel2
rlabel metal1 -783 226 -783 226 1 CLK
rlabel metal1 -780 202 -780 202 1 Imm0
rlabel metal1 -780 194 -780 194 1 Imm1
rlabel metal1 -780 186 -780 186 1 Imm2
rlabel metal1 -780 178 -780 178 1 Imm3
rlabel metal1 -780 170 -780 170 1 Imm4
rlabel metal1 -780 162 -780 162 1 Imm5
rlabel metal1 -780 154 -780 154 1 Imm6
rlabel metal1 -780 146 -780 146 1 Imm7
rlabel metal1 -782 242 -782 242 1 Imm_en
rlabel metal2 -547 342 -547 342 5 C0
rlabel metal2 -483 342 -483 342 5 C1
rlabel metal2 -419 342 -419 342 5 C2
rlabel metal2 -355 341 -355 341 5 C3
rlabel metal2 -291 342 -291 342 5 C4
rlabel metal2 -227 342 -227 342 5 C5
rlabel metal2 -163 342 -163 342 5 C6
rlabel metal2 -99 342 -99 342 5 C7
rlabel metal1 -605 334 -605 334 1 VDD
rlabel metal1 -606 250 -606 250 1 VSS
rlabel metal2 2936 218 2936 218 1 A0
rlabel metal2 2944 218 2944 218 1 A1
rlabel metal2 2952 218 2952 218 1 A2
rlabel metal2 2960 218 2960 218 1 A3
rlabel metal2 2968 218 2968 218 1 A4
rlabel metal2 2976 218 2976 218 1 A5
rlabel metal2 2984 218 2984 218 1 A6
rlabel metal2 2992 218 2992 218 1 A7
rlabel metal2 3000 218 3000 218 1 B0
rlabel metal2 3008 218 3008 218 1 B1
rlabel metal2 3016 218 3016 218 1 B2
rlabel metal2 3024 218 3024 218 1 B3
rlabel metal2 3032 218 3032 218 1 B4
rlabel metal2 3040 218 3040 218 1 B5
rlabel metal2 3048 218 3048 218 1 B6
rlabel metal2 3056 218 3056 218 7 B7
<< end >>
