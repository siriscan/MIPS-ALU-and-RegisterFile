magic
tech scmos
timestamp 1746070328
<< nwell >>
rect 655 738 759 759
rect 655 725 740 738
rect 658 710 686 725
rect 658 343 685 710
rect 654 342 685 343
rect 654 326 689 342
rect 67 311 92 326
rect 684 325 689 326
rect 67 -21 91 311
rect 67 -60 685 -21
rect 658 -328 685 -60
rect 658 -343 686 -328
rect 655 -376 739 -343
rect 954 -362 956 -342
<< metal1 >>
rect 672 743 740 747
rect 0 703 740 707
rect 613 659 740 663
rect 950 636 2014 640
rect 2050 636 2234 640
rect 925 628 2022 632
rect 2058 628 2234 632
rect 900 620 2030 624
rect 2066 620 2234 624
rect 875 612 2038 616
rect 2074 612 2234 616
rect 850 604 2070 608
rect 2082 604 2234 608
rect 825 596 2062 600
rect 2092 596 2234 600
rect 800 587 2054 591
rect 2101 587 2234 591
rect 775 578 2046 582
rect 2109 578 2234 582
rect 2042 570 2078 574
rect 2034 562 2088 566
rect 2026 554 2097 558
rect 2018 546 2105 550
rect 942 505 2063 509
rect 917 497 1872 501
rect 892 489 1682 493
rect 867 481 1493 485
rect 842 473 1305 477
rect 817 464 1114 468
rect 739 455 763 459
rect 792 455 924 459
rect 87 318 134 322
rect 106 234 117 238
rect -29 210 0 214
rect -29 201 0 205
rect -29 193 0 197
rect -29 185 0 189
rect -29 177 0 181
rect -29 169 0 173
rect -29 161 0 165
rect -29 153 0 157
rect 767 -36 2235 -32
rect 87 -42 668 -38
rect 739 -46 763 -42
rect 792 -46 924 -42
rect 928 -46 2235 -42
rect 817 -55 1114 -51
rect 1118 -55 2235 -51
rect 842 -64 1305 -60
rect 1309 -64 2235 -60
rect -2 -69 97 -65
rect 867 -72 1493 -68
rect 1497 -72 2235 -68
rect 892 -80 1682 -76
rect 1686 -80 2235 -76
rect 917 -88 1872 -84
rect 1876 -88 2235 -84
rect 942 -96 2063 -92
rect 2067 -96 2235 -92
rect 647 -135 2235 -131
rect 775 -200 2237 -196
rect 800 -209 2237 -205
rect 825 -218 2237 -214
rect 850 -226 2237 -222
rect 875 -234 2237 -230
rect 900 -242 2237 -238
rect 925 -250 2237 -246
rect 950 -258 2237 -254
rect 613 -281 739 -277
rect 0 -325 740 -321
rect 672 -365 739 -361
<< m2contact >>
rect 668 743 672 747
rect 609 659 613 663
rect 946 636 950 640
rect 2014 636 2018 640
rect 2046 636 2050 640
rect 921 628 925 632
rect 2022 628 2026 632
rect 2054 628 2058 632
rect 896 620 900 624
rect 2030 620 2034 624
rect 2062 620 2066 624
rect 871 612 875 616
rect 2038 612 2042 616
rect 2070 612 2074 616
rect 846 604 850 608
rect 2070 604 2074 608
rect 2078 604 2082 608
rect 821 596 825 600
rect 2062 596 2066 600
rect 2088 596 2092 600
rect 796 587 800 591
rect 2054 587 2058 591
rect 2097 587 2101 591
rect 771 578 775 582
rect 2046 578 2050 582
rect 2105 578 2109 582
rect 2038 570 2042 574
rect 2078 570 2082 574
rect 2030 562 2034 566
rect 2088 562 2092 566
rect 2022 554 2026 558
rect 2097 554 2101 558
rect 2014 546 2018 550
rect 2105 546 2109 550
rect 938 505 942 509
rect 2063 505 2067 509
rect 913 497 917 501
rect 1872 497 1876 501
rect 888 489 892 493
rect 1682 489 1686 493
rect 863 481 867 485
rect 1493 481 1497 485
rect 838 473 842 477
rect 1305 473 1309 477
rect 813 464 817 468
rect 1114 464 1118 468
rect 735 455 739 459
rect 763 455 767 459
rect 788 455 792 459
rect 924 455 928 459
rect 83 318 87 322
rect 668 318 672 322
rect 609 234 613 238
rect 763 -36 767 -32
rect 83 -42 87 -38
rect 668 -42 672 -38
rect 735 -46 739 -42
rect 763 -46 767 -42
rect 788 -46 792 -42
rect 924 -46 928 -42
rect 813 -55 817 -51
rect 1114 -55 1118 -51
rect 838 -64 842 -60
rect 1305 -64 1309 -60
rect 97 -69 101 -65
rect 863 -72 867 -68
rect 1493 -72 1497 -68
rect 888 -80 892 -76
rect 1682 -80 1686 -76
rect 913 -88 917 -84
rect 1872 -88 1876 -84
rect 938 -96 942 -92
rect 2063 -96 2067 -92
rect 643 -135 647 -131
rect 771 -200 775 -196
rect 796 -209 800 -205
rect 821 -218 825 -214
rect 846 -226 850 -222
rect 871 -234 875 -230
rect 896 -242 900 -238
rect 921 -250 925 -246
rect 946 -258 950 -254
rect 609 -281 613 -277
rect 668 -365 672 -361
<< metal2 >>
rect 83 -38 87 318
rect 609 238 613 659
rect 668 322 672 743
rect 763 459 767 703
rect 771 582 775 703
rect 788 459 792 703
rect 796 591 800 703
rect 813 468 817 703
rect 821 600 825 703
rect 838 477 842 703
rect 846 608 850 703
rect 863 485 867 703
rect 871 616 875 703
rect 888 493 892 703
rect 896 624 900 703
rect 913 501 917 703
rect 921 632 925 703
rect 938 509 942 703
rect 946 640 950 703
rect 2014 550 2018 636
rect 2022 558 2026 628
rect 2030 566 2034 620
rect 2038 574 2042 612
rect 2046 582 2050 636
rect 2054 591 2058 628
rect 2062 600 2066 620
rect 2070 608 2074 612
rect 2078 574 2082 604
rect 2088 566 2092 596
rect 2097 558 2101 587
rect 2105 550 2109 578
rect 735 389 739 455
rect 924 381 928 455
rect 1114 373 1118 464
rect 1305 365 1309 473
rect 1493 357 1497 481
rect 1682 349 1686 489
rect 1872 341 1876 497
rect 2063 333 2067 505
rect 97 -65 101 9
rect 609 -277 613 234
rect 643 -131 647 40
rect 668 -361 672 -42
rect 735 -42 739 31
rect 763 -42 767 -36
rect 924 -42 928 27
rect 763 -321 767 -46
rect 771 -321 775 -200
rect 788 -321 792 -46
rect 1114 -51 1118 33
rect 796 -321 800 -209
rect 813 -321 817 -55
rect 1305 -60 1309 33
rect 821 -321 825 -218
rect 838 -321 842 -64
rect 1493 -68 1497 33
rect 846 -321 850 -226
rect 863 -321 867 -72
rect 1682 -76 1686 31
rect 871 -321 875 -234
rect 888 -321 892 -80
rect 1872 -84 1876 33
rect 896 -321 900 -242
rect 913 -321 917 -88
rect 2063 -92 2067 33
rect 921 -321 925 -250
rect 938 -321 942 -96
rect 946 -321 950 -258
use BUFFER8  BUFFER8_0
timestamp 1746041965
transform 1 0 738 0 -1 -277
box -4 -8 218 91
use BUFFER8  BUFFER8_1
timestamp 1746041965
transform 1 0 738 0 1 659
box -4 -8 218 91
use reg8_8bitMUX2to1  reg8_8bitMUX2to1_0
timestamp 1746070328
transform 1 0 91 0 1 218
box -91 -218 2032 171
<< labels >>
rlabel metal1 -27 212 -27 212 1 C0
rlabel metal1 -27 203 -27 203 1 C1
rlabel metal1 -27 195 -27 195 1 C2
rlabel metal1 -27 187 -27 187 1 C3
rlabel metal1 -27 179 -27 179 1 C4
rlabel metal1 -27 171 -27 171 1 C5
rlabel metal1 -27 163 -27 163 1 C6
rlabel metal1 -27 155 -27 155 1 C7
rlabel metal1 2 705 2 705 1 b_en
rlabel metal1 125 320 125 320 1 VDD
rlabel metal1 111 236 111 236 1 VSS
rlabel metal1 0 -67 0 -67 1 reg_en
rlabel metal1 2232 638 2232 638 1 B0
rlabel metal1 2232 630 2232 630 1 B1
rlabel metal1 2232 622 2232 622 1 B2
rlabel metal1 2232 614 2232 614 1 B3
rlabel metal1 2232 606 2232 606 1 B4
rlabel metal1 2232 598 2232 598 1 B5
rlabel metal1 2232 589 2232 589 1 B6
rlabel metal1 2232 580 2232 580 1 B7
rlabel metal1 2233 -34 2233 -34 1 Q0
rlabel metal1 2233 -44 2233 -44 1 Q1
rlabel metal1 2233 -53 2233 -53 1 Q2
rlabel metal1 2233 -62 2233 -62 1 Q3
rlabel metal1 2233 -70 2233 -70 1 Q4
rlabel metal1 2233 -78 2233 -78 1 Q5
rlabel metal1 2233 -86 2233 -86 1 Q6
rlabel metal1 2233 -94 2233 -94 1 Q7
rlabel metal1 2233 -133 2233 -133 1 CLK
rlabel metal1 2 -323 2 -323 1 a_en
rlabel metal1 2235 -256 2235 -256 1 A7
rlabel metal1 2235 -248 2235 -248 1 A6
rlabel metal1 2235 -240 2235 -240 1 A5
rlabel metal1 2235 -232 2235 -232 1 A4
rlabel metal1 2235 -224 2235 -224 1 A3
rlabel metal1 2235 -216 2235 -216 1 A2
rlabel metal1 2235 -207 2235 -207 1 A1
rlabel metal1 2235 -198 2235 -198 1 A0
<< end >>
