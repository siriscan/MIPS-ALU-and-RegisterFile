magic
tech scmos
timestamp 1746041965
<< polycontact >>
rect 16 37 20 41
rect 56 37 60 41
rect 96 37 100 41
rect 136 37 140 41
rect 176 37 180 41
rect 216 37 220 41
rect 256 37 260 41
rect 296 37 300 41
rect 8 23 12 27
rect 48 23 52 27
rect 88 23 92 27
rect 128 23 132 27
rect 168 23 172 27
rect 208 23 212 27
rect 248 23 252 27
rect 288 23 292 27
<< metal1 >>
rect 5 84 15 88
rect 39 26 43 30
rect 79 27 83 31
rect 119 26 123 30
rect 159 26 163 30
rect 199 25 203 29
rect 239 27 243 31
rect 279 28 283 32
rect 319 28 323 32
rect 5 0 13 4
use AND2  AND2_7
timestamp 1740126148
transform 1 0 285 0 1 0
box -5 0 45 92
use AND2  AND2_6
timestamp 1740126148
transform 1 0 245 0 1 0
box -5 0 45 92
use AND2  AND2_5
timestamp 1740126148
transform 1 0 205 0 1 0
box -5 0 45 92
use AND2  AND2_4
timestamp 1740126148
transform 1 0 165 0 1 0
box -5 0 45 92
use AND2  AND2_3
timestamp 1740126148
transform 1 0 125 0 1 0
box -5 0 45 92
use AND2  AND2_2
timestamp 1740126148
transform 1 0 85 0 1 0
box -5 0 45 92
use AND2  AND2_1
timestamp 1740126148
transform 1 0 45 0 1 0
box -5 0 45 92
use AND2  AND2_0
timestamp 1740126148
transform 1 0 5 0 1 0
box -5 0 45 92
<< labels >>
rlabel metal1 9 86 9 86 1 VDD
rlabel metal1 9 2 9 2 1 VSS
rlabel polycontact 10 25 10 25 1 A0
rlabel polycontact 50 25 50 25 1 A1
rlabel polycontact 90 25 90 25 1 A2
rlabel polycontact 130 25 130 25 1 A3
rlabel polycontact 170 25 170 25 1 A4
rlabel polycontact 210 25 210 25 1 A5
rlabel polycontact 250 25 250 25 1 A6
rlabel polycontact 290 25 290 25 1 A7
rlabel polycontact 18 39 18 39 1 B0
rlabel polycontact 58 39 58 39 1 B1
rlabel polycontact 98 39 98 39 1 B2
rlabel polycontact 138 39 138 39 1 B3
rlabel polycontact 178 39 178 39 1 B4
rlabel polycontact 218 39 218 39 1 B5
rlabel polycontact 258 39 258 39 1 B6
rlabel polycontact 298 39 298 39 1 B7
rlabel metal1 41 28 41 28 1 Y0
rlabel metal1 81 29 81 29 1 Y1
rlabel metal1 121 28 121 28 1 Y2
rlabel metal1 161 28 161 28 1 Y3
rlabel metal1 201 27 201 27 1 Y4
rlabel metal1 241 29 241 29 1 Y5
rlabel metal1 281 30 281 30 1 Y6
rlabel metal1 321 30 321 30 1 Y7
<< end >>
