magic
tech scmos
timestamp 1742676329
<< metal1 >>
rect 0 0 4 88
<< end >>
