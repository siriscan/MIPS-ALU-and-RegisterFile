magic
tech scmos
timestamp 1741159115
<< nwell >>
rect -4 32 36 91
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
rect 23 8 25 12
<< ptransistor >>
rect 7 38 9 42
rect 15 38 17 42
rect 23 38 25 42
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
rect 14 8 15 12
rect 17 8 23 12
rect 25 8 26 12
<< pdiffusion >>
rect 6 38 7 42
rect 9 38 10 42
rect 14 38 15 42
rect 17 38 18 42
rect 22 38 23 42
rect 25 38 26 42
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
rect 26 8 30 12
<< pdcontact >>
rect 2 38 6 42
rect 10 38 14 42
rect 18 38 22 42
rect 26 38 30 42
<< psubstratepcontact >>
rect 2 0 6 4
rect 26 0 30 4
<< nsubstratencontact >>
rect 2 84 6 88
<< polysilicon >>
rect 7 42 9 44
rect 15 42 17 44
rect 23 42 25 44
rect 7 37 9 38
rect 5 35 9 37
rect 5 25 7 35
rect 5 23 9 25
rect 7 20 9 23
rect 6 16 9 20
rect 7 12 9 16
rect 15 12 17 38
rect 23 20 25 38
rect 23 16 26 20
rect 23 12 25 16
rect 7 6 9 8
rect 15 6 17 8
rect 23 6 25 8
<< polycontact >>
rect 11 28 15 32
rect 2 16 6 20
rect 26 16 30 20
<< metal1 >>
rect 0 84 2 88
rect 6 84 32 88
rect 2 42 6 84
rect 10 45 30 49
rect 10 42 14 45
rect 26 42 30 45
rect 18 20 22 38
rect 10 16 22 20
rect 10 12 14 16
rect 2 4 6 8
rect 26 4 30 8
rect 0 0 2 4
rect 6 0 26 4
rect 30 0 32 4
<< labels >>
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel psubstratepcontact 28 2 28 2 1 VSS
rlabel polycontact 4 18 4 18 1 A
rlabel polycontact 13 30 13 30 1 B
rlabel polycontact 28 18 28 18 1 C
rlabel metal1 20 24 20 24 1 Y
rlabel nsubstratencontact 4 86 4 86 1 VDD
<< end >>
