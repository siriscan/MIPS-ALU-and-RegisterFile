magic
tech scmos
timestamp 1746597901
<< nwell >>
rect 2039 252 2043 256
<< metal1 >>
rect 8 252 12 256
rect 2039 252 2484 256
rect 9 168 13 172
rect 2038 168 2484 172
rect 8 160 12 164
rect 8 144 12 148
rect -6 120 1 124
rect 2104 120 2924 124
rect -6 112 1 116
rect 2100 112 2151 116
rect 2155 112 2924 116
rect -6 104 1 108
rect 2100 104 2202 108
rect 2206 104 2924 108
rect -6 96 1 100
rect 2100 96 2253 100
rect 2257 96 2924 100
rect -6 88 1 92
rect 2100 88 2304 92
rect 2308 88 2924 92
rect -6 80 1 84
rect 2100 80 2355 84
rect 2359 80 2924 84
rect -6 72 1 76
rect 2100 72 2406 76
rect 2410 72 2924 76
rect -6 64 1 68
rect 2100 64 2457 68
rect 2461 64 2924 68
rect 2050 56 2063 60
rect 2067 56 2490 60
rect 2494 56 2924 60
rect 2050 48 2114 52
rect 2118 48 2541 52
rect 2545 48 2924 52
rect 2050 40 2165 44
rect 2169 40 2592 44
rect 2596 40 2924 44
rect 2050 32 2216 36
rect 2220 32 2643 36
rect 2647 32 2924 36
rect 2050 24 2267 28
rect 2271 24 2694 28
rect 2698 24 2924 28
rect 2050 16 2318 20
rect 2322 16 2745 20
rect 2749 16 2924 20
rect 2050 8 2369 12
rect 2373 8 2796 12
rect 2800 8 2924 12
rect 2050 0 2420 4
rect 2424 0 2847 4
rect 2851 0 2924 4
rect 2531 -8 2924 -4
rect 2527 -16 2578 -12
rect 2582 -16 2924 -12
rect 2527 -24 2629 -20
rect 2633 -24 2924 -20
rect 2527 -32 2680 -28
rect 2684 -32 2924 -28
rect 2527 -40 2731 -36
rect 2735 -40 2924 -36
rect 2527 -48 2782 -44
rect 2786 -48 2924 -44
rect 0 -56 2047 -52
rect 2527 -56 2833 -52
rect 2837 -56 2924 -52
rect 0 -64 2474 -60
rect 2527 -64 2884 -60
rect 2888 -64 2924 -60
<< m2contact >>
rect 2100 120 2104 124
rect 2151 112 2155 116
rect 2202 104 2206 108
rect 2253 96 2257 100
rect 2304 88 2308 92
rect 2355 80 2359 84
rect 2406 72 2410 76
rect 2457 64 2461 68
rect 2063 56 2067 60
rect 2490 56 2494 60
rect 2114 48 2118 52
rect 2541 48 2545 52
rect 2165 40 2169 44
rect 2592 40 2596 44
rect 2216 32 2220 36
rect 2643 32 2647 36
rect 2267 24 2271 28
rect 2694 24 2698 28
rect 2318 16 2322 20
rect 2745 16 2749 20
rect 2369 8 2373 12
rect 2796 8 2800 12
rect 2420 0 2424 4
rect 2847 0 2851 4
rect 2527 -8 2531 -4
rect 2578 -16 2582 -12
rect 2629 -24 2633 -20
rect 2680 -32 2684 -28
rect 2731 -40 2735 -36
rect 2782 -48 2786 -44
rect 2047 -56 2051 -52
rect 2833 -56 2837 -52
rect 2474 -64 2478 -60
rect 2884 -64 2888 -60
<< metal2 >>
rect 2047 -52 2051 212
rect 2063 60 2067 156
rect 2100 124 2104 156
rect 2114 52 2118 156
rect 2151 116 2155 156
rect 2165 44 2169 156
rect 2202 108 2206 156
rect 2216 36 2220 156
rect 2253 100 2257 156
rect 2267 28 2271 156
rect 2304 92 2308 156
rect 2318 20 2322 156
rect 2355 84 2359 156
rect 2369 12 2373 156
rect 2406 76 2410 156
rect 2420 4 2424 156
rect 2457 68 2461 156
rect 2474 -60 2478 212
rect 2490 60 2494 156
rect 2527 -4 2531 156
rect 2541 52 2545 156
rect 2578 -12 2582 156
rect 2592 44 2596 156
rect 2629 -20 2633 156
rect 2643 36 2647 156
rect 2680 -28 2684 156
rect 2694 28 2698 156
rect 2731 -36 2735 156
rect 2745 20 2749 156
rect 2782 -44 2786 156
rect 2796 12 2800 156
rect 2833 -52 2837 156
rect 2847 4 2851 156
rect 2884 -60 2888 156
use REGv2  REGv2_0
timestamp 1746512792
transform 1 0 531 0 1 120
box -531 -120 1519 140
use BUFFER8v2  BUFFER8v2_1
timestamp 1746552068
transform 1 0 2468 0 1 160
box -3 -4 444 104
use BUFFER8v2  BUFFER8v2_0
timestamp 1746552068
transform 1 0 2041 0 1 160
box -3 -4 444 104
<< labels >>
rlabel metal1 10 146 10 146 1 CLK
rlabel metal1 10 162 10 162 1 reg_en
rlabel metal1 11 170 11 170 1 VSS
rlabel metal1 10 254 10 254 1 VDD
rlabel metal1 -4 122 -4 122 3 C0
rlabel metal1 -4 114 -4 114 3 C1
rlabel metal1 -4 106 -4 106 3 C2
rlabel metal1 -4 98 -4 98 3 C3
rlabel metal1 -4 90 -4 90 3 C4
rlabel metal1 -4 82 -4 82 3 C5
rlabel metal1 -4 74 -4 74 3 C6
rlabel metal1 -4 66 -4 66 3 C7
rlabel metal1 2921 2 2921 2 8 Q7
rlabel metal1 2922 10 2922 10 7 Q6
rlabel metal1 2921 18 2921 18 7 Q5
rlabel metal1 2921 26 2921 26 7 Q4
rlabel metal1 2921 34 2921 34 7 Q3
rlabel metal1 2921 42 2921 42 7 Q2
rlabel metal1 2922 50 2922 50 7 Q1
rlabel metal1 2922 58 2922 58 7 Q0
rlabel metal1 2914 -6 2914 -6 7 B0
rlabel metal1 2914 -14 2914 -14 7 B1
rlabel metal1 2914 -22 2914 -22 7 B2
rlabel metal1 2914 -30 2914 -30 7 B3
rlabel metal1 2914 -38 2914 -38 7 B4
rlabel metal1 2913 -46 2913 -46 7 B5
rlabel metal1 2914 -54 2914 -54 7 B6
rlabel metal1 2914 -62 2914 -62 8 B7
rlabel metal1 2923 122 2923 122 7 A0
rlabel metal1 2922 114 2922 114 7 A1
rlabel metal1 2923 106 2923 106 7 A2
rlabel metal1 2922 98 2922 98 7 A3
rlabel metal1 2922 90 2922 90 7 A4
rlabel metal1 2922 82 2922 82 7 A5
rlabel metal1 2921 74 2921 74 7 A6
rlabel metal1 2922 66 2922 66 7 A7
rlabel metal1 3 -54 3 -54 2 a_enb
rlabel metal1 3 -62 3 -62 2 b_enb
<< end >>
