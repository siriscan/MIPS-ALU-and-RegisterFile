magic
tech scmos
timestamp 1741221840
<< metal1 >>
rect 5 84 9 88
rect 25 58 29 62
rect 17 41 21 45
rect 40 29 44 40
rect 48 34 52 52
rect 8 24 12 28
rect 36 25 44 29
rect 17 0 21 4
use INV  INV_0
timestamp 1741159900
transform 1 0 38 0 1 0
box -4 0 20 91
use NAND3  NAND3_0
timestamp 1741221395
transform 1 0 5 0 1 0
box -5 0 38 91
<< labels >>
rlabel metal1 7 86 7 86 1 VDD
rlabel metal1 27 60 27 60 1 C
rlabel metal1 19 43 19 43 1 B
rlabel metal1 10 26 10 26 1 A
rlabel metal1 19 2 19 2 1 VSS
rlabel metal1 50 44 50 44 1 Y
<< end >>
