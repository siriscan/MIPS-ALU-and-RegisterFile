magic
tech scmos
timestamp 1746652338
<< metal1 >>
rect 246 2681 7951 2685
rect 310 2673 7959 2677
rect 374 2665 7967 2669
rect 438 2657 7975 2661
rect 502 2649 7983 2653
rect 566 2641 7991 2645
rect 630 2633 7999 2637
rect 694 2625 8007 2629
rect 178 2608 183 2612
rect 178 2524 183 2528
rect 2 2516 6 2520
rect 2 2500 6 2504
rect 2 2476 6 2480
rect 2 2468 6 2472
rect 2 2460 6 2464
rect 2 2452 6 2456
rect 8011 2451 8015 2455
rect 2 2444 6 2448
rect 8011 2443 8015 2447
rect 2 2436 6 2440
rect 8011 2435 8015 2439
rect 2 2428 6 2432
rect 8011 2427 8015 2431
rect 2 2420 6 2424
rect 8011 2419 8015 2423
rect 3706 2412 3711 2416
rect 3729 2412 3849 2416
rect 3854 2412 3858 2416
rect 8011 2411 8015 2415
rect 3706 2404 3711 2408
rect 3737 2404 3849 2408
rect 3854 2404 3858 2408
rect 8011 2403 8015 2407
rect 3706 2396 3711 2400
rect 3745 2396 3849 2400
rect 3854 2396 3858 2400
rect 8011 2395 8015 2399
rect 3706 2388 3711 2392
rect 3753 2388 3849 2392
rect 3854 2388 3858 2392
rect 8011 2387 8015 2391
rect 3706 2380 3711 2384
rect 3761 2380 3849 2384
rect 3854 2380 3858 2384
rect 3706 2372 3711 2376
rect 3769 2372 3849 2376
rect 3854 2372 3858 2376
rect 3706 2364 3711 2368
rect 3777 2364 3849 2368
rect 3854 2364 3858 2368
rect 3706 2356 3711 2360
rect 3785 2356 3849 2360
rect 3854 2356 3858 2360
rect 3854 2348 3858 2352
rect 3854 2340 3858 2344
rect 3854 2332 3858 2336
rect 3854 2324 3858 2328
rect 3854 2316 3858 2320
rect 3854 2308 3858 2312
rect 3854 2300 3858 2304
rect 3854 2292 3858 2296
rect 12 2176 26 2180
rect 12 2168 26 2172
rect 12 2152 26 2156
rect 12 2136 26 2140
rect 3709 2072 3713 2076
rect 3709 2064 3713 2068
rect 3709 2056 3713 2060
rect 3709 2048 3713 2052
rect 3709 2040 3713 2044
rect 3709 2032 3713 2036
rect 3709 2024 3713 2028
rect 3709 2016 3713 2020
rect 12 1933 26 1937
rect 12 1917 26 1921
rect 12 1901 26 1905
rect 3709 1732 3713 1736
rect 3709 1724 3713 1728
rect 3709 1716 3713 1720
rect 3709 1708 3713 1712
rect 3709 1700 3713 1704
rect 3709 1692 3713 1696
rect 11 1685 22 1689
rect 3709 1684 3713 1688
rect 3709 1676 3713 1680
rect 11 1669 22 1673
rect 11 1653 22 1657
rect 3708 1392 3712 1396
rect 3708 1384 3712 1388
rect 3708 1376 3712 1380
rect 3708 1368 3712 1372
rect 3708 1360 3712 1364
rect 3708 1352 3712 1356
rect 3708 1344 3712 1348
rect 3708 1336 3712 1340
rect 3710 1052 3714 1056
rect 3710 1044 3714 1048
rect 3710 1036 3714 1040
rect 3710 1028 3714 1032
rect 3710 1020 3714 1024
rect 3710 1012 3714 1016
rect 3710 1004 3714 1008
rect 3710 996 3714 1000
rect 3709 712 3713 716
rect 3709 704 3713 708
rect 3709 696 3713 700
rect 3709 688 3713 692
rect 3709 680 3713 684
rect 3709 672 3713 676
rect 3709 664 3713 668
rect 3709 656 3713 660
rect 3707 372 3711 376
rect 3707 364 3711 368
rect 3707 356 3711 360
rect 3707 348 3711 352
rect 3707 340 3711 344
rect 3707 332 3711 336
rect 3707 324 3711 328
rect 3707 316 3711 320
rect 613 136 642 140
<< m2contact >>
rect 242 2681 246 2685
rect 7951 2681 7955 2685
rect 306 2673 310 2677
rect 7959 2673 7963 2677
rect 370 2665 374 2669
rect 7967 2665 7971 2669
rect 434 2657 438 2661
rect 7975 2657 7979 2661
rect 498 2649 502 2653
rect 7983 2649 7987 2653
rect 562 2641 566 2645
rect 7991 2641 7995 2645
rect 626 2633 630 2637
rect 7999 2633 8003 2637
rect 690 2625 694 2629
rect 8007 2625 8011 2629
rect 3696 2608 3700 2612
rect 3701 2524 3705 2528
rect 3899 2476 3903 2480
rect 3879 2467 3883 2471
rect 3912 2459 3916 2463
rect 3920 2451 3924 2455
rect 3928 2443 3932 2447
rect 3725 2412 3729 2416
rect 3733 2404 3737 2408
rect 3741 2396 3745 2400
rect 3749 2388 3753 2392
rect 3757 2380 3761 2384
rect 3765 2372 3769 2376
rect 3773 2364 3777 2368
rect 3781 2356 3785 2360
rect 3876 1259 3880 1263
rect 3853 1171 3857 1175
<< metal2 >>
rect 242 2619 246 2681
rect 306 2620 310 2673
rect 370 2619 374 2665
rect 434 2618 438 2657
rect 498 2619 502 2649
rect 562 2620 566 2641
rect 626 2620 630 2633
rect 690 2617 694 2625
rect 3912 2463 3916 2700
rect 3920 2455 3924 2700
rect 3928 2447 3932 2700
rect 7951 2426 7955 2681
rect 7959 2426 7963 2673
rect 7967 2426 7971 2665
rect 7975 2421 7979 2657
rect 3725 2356 3729 2412
rect 3733 2408 3737 2416
rect 3733 2356 3737 2404
rect 3741 2400 3745 2416
rect 3741 2356 3745 2396
rect 3749 2392 3753 2416
rect 3749 2356 3753 2388
rect 3757 2384 3761 2416
rect 3757 2356 3761 2380
rect 3765 2376 3769 2416
rect 3765 2356 3769 2372
rect 3773 2368 3777 2416
rect 3773 2356 3777 2364
rect 3781 2360 3785 2416
rect 7983 2394 7987 2649
rect 7991 2399 7995 2641
rect 7999 2392 8003 2633
rect 8007 2391 8011 2625
rect 3853 -12 3857 1171
rect 3876 -12 3880 1259
<< m3contact >>
rect 3700 2608 3704 2612
rect 3705 2524 3709 2528
rect 3903 2476 3907 2480
rect 3879 2471 3883 2475
<< metal3 >>
rect 3699 2612 3908 2613
rect 3699 2608 3700 2612
rect 3704 2608 3908 2612
rect 3699 2607 3908 2608
rect 3704 2528 3885 2529
rect 3704 2524 3705 2528
rect 3709 2524 3885 2528
rect 3704 2523 3885 2524
rect 3878 2475 3885 2523
rect 3902 2480 3908 2607
rect 3902 2476 3903 2480
rect 3907 2476 3908 2480
rect 3902 2475 3908 2476
rect 3878 2471 3879 2475
rect 3883 2471 3885 2475
rect 3878 2470 3885 2471
use REGISTER_FILEv2  REGISTER_FILEv2_0
timestamp 1746652306
transform 1 0 791 0 1 2276
box -791 -2276 3058 345
use ALU  ALU_0
timestamp 1746489366
transform 1 0 4266 0 1 767
box -417 0 3745 1796
<< labels >>
rlabel metal1 180 2526 180 2526 1 VSS
rlabel metal1 181 2610 181 2610 1 VDD
rlabel metal1 3855 2414 3855 2414 3 A0
rlabel metal1 3855 2406 3855 2406 3 A1
rlabel metal1 3855 2398 3855 2398 3 A2
rlabel metal1 3855 2390 3855 2390 3 A3
rlabel metal1 3855 2382 3855 2382 3 A4
rlabel metal1 3855 2374 3855 2374 3 A5
rlabel metal1 3855 2366 3855 2366 3 A6
rlabel metal1 3855 2358 3855 2358 3 A7
rlabel metal1 3855 2350 3855 2350 3 B0
rlabel metal1 3855 2342 3855 2342 3 B1
rlabel metal1 3855 2334 3855 2334 3 B2
rlabel metal1 3855 2326 3855 2326 3 B3
rlabel metal1 3855 2318 3855 2318 3 B4
rlabel metal1 3855 2310 3855 2310 3 B5
rlabel metal1 3855 2302 3855 2302 3 B6
rlabel metal1 3855 2294 3855 2294 3 B7
rlabel metal2 3914 2698 3914 2698 5 func0
rlabel metal2 3922 2698 3922 2698 5 func1
rlabel metal2 3930 2698 3930 2698 5 func2
rlabel metal1 4 2518 4 2518 3 imm_en
rlabel metal1 4 2478 4 2478 1 Imm0
rlabel metal1 4 2470 4 2470 1 Imm1
rlabel metal1 4 2462 4 2462 1 Imm2
rlabel metal1 4 2454 4 2454 1 Imm3
rlabel metal1 4 2446 4 2446 1 Imm4
rlabel metal1 4 2438 4 2438 1 Imm5
rlabel metal1 4 2430 4 2430 1 Imm6
rlabel metal1 4 2422 4 2422 1 Imm7
rlabel space 10 3855 10 3855 5 RorL
rlabel metal2 3855 -10 3855 -10 1 RorL
rlabel metal2 3878 -10 3878 -10 1 LorA
rlabel metal1 17 2178 17 2178 1 Write_Address3
rlabel metal1 17 2170 17 2170 1 Write_Address0
rlabel metal1 17 2154 17 2154 1 Write_Address1
rlabel metal1 17 2138 17 2138 1 Write_Address2
rlabel metal1 17 1935 17 1935 1 A_Read_Address0
rlabel metal1 17 1919 17 1919 1 A_Read_Address1
rlabel metal1 17 1903 17 1903 1 A_Read_Address2
rlabel metal1 14 1687 14 1687 1 B_Read_Address0
rlabel metal1 14 1671 14 1671 1 B_Read_Address1
rlabel metal1 14 1655 14 1655 1 B_Read_Address2
rlabel metal1 4 2502 4 2502 3 clk
rlabel metal1 3708 2414 3708 2414 1 reg_zero0
rlabel metal1 3708 2406 3708 2406 1 reg_zero1
rlabel metal1 3708 2398 3708 2398 1 reg_zero2
rlabel metal1 3708 2390 3708 2390 1 reg_zero3
rlabel metal1 3708 2382 3708 2382 1 reg_zero4
rlabel metal1 3708 2374 3708 2374 1 reg_zero5
rlabel metal1 3708 2366 3708 2366 1 reg_zero6
rlabel metal1 3708 2358 3708 2358 1 reg_zero7
rlabel metal1 3712 2074 3712 2074 1 reg_one0
rlabel metal1 3712 2066 3712 2066 1 reg_one1
rlabel metal1 3712 2058 3712 2058 1 reg_one2
rlabel metal1 3712 2050 3712 2050 1 reg_one3
rlabel metal1 3712 2042 3712 2042 1 reg_one4
rlabel metal1 3712 2034 3712 2034 1 reg_one5
rlabel metal1 3712 2026 3712 2026 1 reg_one6
rlabel metal1 3712 2018 3712 2018 1 reg_one7
rlabel metal1 3712 1734 3712 1734 1 reg_two0
rlabel metal1 3712 1726 3712 1726 1 reg_two1
rlabel metal1 3712 1718 3712 1718 1 reg_two2
rlabel metal1 3712 1710 3712 1710 1 reg_two3
rlabel metal1 3711 1702 3711 1702 1 reg_two4
rlabel metal1 3712 1694 3712 1694 1 reg_two5
rlabel metal1 3712 1686 3712 1686 1 reg_two6
rlabel metal1 3712 1678 3712 1678 1 reg_two7
rlabel metal1 3711 1394 3711 1394 1 reg_three0
rlabel metal1 3711 1386 3711 1386 1 reg_three1
rlabel metal1 3711 1378 3711 1378 1 reg_three2
rlabel metal1 3711 1370 3711 1370 1 reg_three3
rlabel metal1 3711 1362 3711 1362 1 reg_three4
rlabel metal1 3711 1354 3711 1354 1 reg_three5
rlabel metal1 3711 1346 3711 1346 1 reg_three6
rlabel metal1 3711 1338 3711 1338 1 reg_three7
rlabel metal1 3713 1054 3713 1054 1 reg_four0
rlabel metal1 3713 1046 3713 1046 1 reg_four1
rlabel metal1 3713 1038 3713 1038 1 reg_four2
rlabel metal1 3713 1030 3713 1030 1 reg_four3
rlabel metal1 3713 1022 3713 1022 1 reg_four4
rlabel metal1 3713 1014 3713 1014 1 reg_four5
rlabel metal1 3714 1006 3714 1006 1 reg_four6
rlabel metal1 3714 998 3714 998 1 reg_four7
rlabel metal1 3713 714 3713 714 1 reg_five0
rlabel metal1 3713 706 3713 706 1 reg_five1
rlabel metal1 3712 698 3712 698 1 reg_five2
rlabel metal1 3712 690 3712 690 1 reg_five3
rlabel metal1 3712 682 3712 682 1 reg_five4
rlabel metal1 3712 674 3712 674 1 reg_five5
rlabel metal1 3712 666 3712 666 1 reg_five6
rlabel metal1 3712 658 3712 658 1 reg_five7
rlabel metal1 3710 374 3710 374 1 reg_six0
rlabel metal1 3710 366 3710 366 1 reg_six1
rlabel metal1 3710 358 3710 358 1 reg_six2
rlabel metal1 3710 350 3710 350 1 reg_six3
rlabel metal1 3710 342 3710 342 1 reg_six4
rlabel metal1 3710 334 3710 334 1 reg_six5
rlabel metal1 3710 326 3710 326 1 reg_six6
rlabel metal1 3710 318 3710 318 1 reg_six7
rlabel metal1 8013 2445 8013 2445 7 Y0
rlabel metal1 8012 2437 8012 2437 7 Y1
rlabel metal1 8012 2429 8012 2429 7 Y2
rlabel metal1 8011 2421 8011 2421 7 Y3
rlabel metal1 8012 2413 8012 2413 7 Y4
rlabel metal1 8012 2405 8012 2405 7 Y5
rlabel metal1 8012 2397 8012 2397 7 Y6
rlabel metal1 8013 2389 8013 2389 7 Y7
rlabel metal1 8012 2453 8012 2453 7 Overflow
<< end >>
