magic
tech scmos
timestamp 1741246353
<< nwell >>
rect -4 69 45 91
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
rect 23 8 25 12
rect 32 8 34 12
<< ptransistor >>
rect 7 76 9 80
rect 15 76 17 80
rect 23 76 25 80
rect 32 76 34 80
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
rect 14 8 15 12
rect 17 8 18 12
rect 22 8 23 12
rect 25 8 27 12
rect 31 8 32 12
rect 34 8 35 12
<< pdiffusion >>
rect 6 76 7 80
rect 9 76 15 80
rect 17 76 23 80
rect 25 76 32 80
rect 34 76 35 80
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
rect 18 8 22 12
rect 27 8 31 12
rect 35 8 39 12
<< pdcontact >>
rect 2 76 6 80
rect 35 76 39 80
<< psubstratepcontact >>
rect 10 0 14 4
rect 27 0 31 4
<< nsubstratencontact >>
rect 2 84 6 88
<< polysilicon >>
rect 7 80 9 82
rect 15 80 17 82
rect 23 80 25 82
rect 32 80 34 82
rect 7 30 9 76
rect 15 40 17 76
rect 23 49 25 76
rect 24 45 25 49
rect 16 36 17 40
rect 8 26 9 30
rect 7 12 9 26
rect 15 12 17 36
rect 23 12 25 45
rect 32 12 34 76
rect 7 6 9 8
rect 15 6 17 8
rect 23 6 25 8
rect 32 6 34 8
<< polycontact >>
rect 28 56 32 60
rect 20 45 24 49
rect 12 36 16 40
rect 4 26 8 30
<< metal1 >>
rect 0 84 2 88
rect 6 84 41 88
rect 2 80 6 84
rect 35 20 39 76
rect 2 16 39 20
rect 2 12 6 16
rect 18 12 22 16
rect 35 12 39 16
rect 10 4 14 8
rect 27 4 31 8
rect 0 0 10 4
rect 14 0 27 4
rect 31 0 41 4
<< labels >>
rlabel psubstratepcontact 12 2 12 2 1 VSS
rlabel psubstratepcontact 29 2 29 2 1 VSS
rlabel polycontact 6 28 6 28 1 A
rlabel polycontact 14 38 14 38 1 B
rlabel polycontact 22 47 22 47 1 C
rlabel polycontact 30 58 30 58 1 D
rlabel metal1 37 42 37 42 1 Y
rlabel nsubstratencontact 4 86 4 86 1 VDD
<< end >>
