magic
tech scmos
timestamp 1746042099
<< nwell >>
rect 685 669 788 696
rect 688 654 716 669
rect 688 39 715 654
rect 688 24 716 39
rect 685 -2 788 24
<< metal1 >>
rect 702 687 768 691
rect 30 647 770 651
rect 643 603 769 607
rect 980 580 2044 584
rect 2080 580 2264 584
rect 955 572 2052 576
rect 2088 572 2264 576
rect 930 564 2060 568
rect 2096 564 2264 568
rect 905 556 2068 560
rect 2104 556 2264 560
rect 880 548 2100 552
rect 2112 548 2264 552
rect 855 540 2092 544
rect 2122 540 2264 544
rect 830 531 2084 535
rect 2131 531 2264 535
rect 805 522 2076 526
rect 2139 522 2264 526
rect 2072 514 2108 518
rect 2064 506 2118 510
rect 2056 498 2127 502
rect 2048 490 2135 494
rect 972 449 2093 453
rect 947 441 1902 445
rect 922 433 1712 437
rect 897 425 1523 429
rect 872 417 1335 421
rect 847 408 1144 412
rect 769 399 793 403
rect 822 399 954 403
rect 643 368 765 372
rect 769 368 954 372
rect 958 368 1144 372
rect 1148 368 1335 372
rect 1339 368 1523 372
rect 1527 368 1712 372
rect 1716 368 1902 372
rect 1906 368 2093 372
rect 797 331 2265 335
rect 769 321 793 325
rect 822 321 954 325
rect 958 321 2265 325
rect 847 312 1144 316
rect 1148 312 2265 316
rect 872 303 1335 307
rect 1339 303 2265 307
rect 897 295 1523 299
rect 1527 295 2265 299
rect 922 287 1712 291
rect 1716 287 2265 291
rect 947 279 1902 283
rect 1906 279 2265 283
rect 972 271 2093 275
rect 2097 271 2265 275
rect 805 167 2267 171
rect 830 158 2267 162
rect 855 149 2267 153
rect 880 141 2267 145
rect 905 133 2267 137
rect 930 125 2267 129
rect 955 117 2267 121
rect 980 109 2267 113
rect 643 86 769 90
rect 30 42 770 46
rect 702 2 770 6
<< m2contact >>
rect 698 687 702 691
rect 639 603 643 607
rect 976 580 980 584
rect 2044 580 2048 584
rect 2076 580 2080 584
rect 951 572 955 576
rect 2052 572 2056 576
rect 2084 572 2088 576
rect 926 564 930 568
rect 2060 564 2064 568
rect 2092 564 2096 568
rect 901 556 905 560
rect 2068 556 2072 560
rect 2100 556 2104 560
rect 876 548 880 552
rect 2100 548 2104 552
rect 2108 548 2112 552
rect 851 540 855 544
rect 2092 540 2096 544
rect 2118 540 2122 544
rect 826 531 830 535
rect 2084 531 2088 535
rect 2127 531 2131 535
rect 801 522 805 526
rect 2076 522 2080 526
rect 2135 522 2139 526
rect 2068 514 2072 518
rect 2108 514 2112 518
rect 2060 506 2064 510
rect 2118 506 2122 510
rect 2052 498 2056 502
rect 2127 498 2131 502
rect 2044 490 2048 494
rect 2135 490 2139 494
rect 968 449 972 453
rect 2093 449 2097 453
rect 943 441 947 445
rect 1902 441 1906 445
rect 918 433 922 437
rect 1712 433 1716 437
rect 893 425 897 429
rect 1523 425 1527 429
rect 868 417 872 421
rect 1335 417 1339 421
rect 843 408 847 412
rect 1144 408 1148 412
rect 765 399 769 403
rect 793 399 797 403
rect 818 399 822 403
rect 954 399 958 403
rect 639 368 643 372
rect 765 368 769 372
rect 954 368 958 372
rect 1144 368 1148 372
rect 1335 368 1339 372
rect 1523 368 1527 372
rect 1712 368 1716 372
rect 1902 368 1906 372
rect 2093 368 2097 372
rect 793 331 797 335
rect 765 321 769 325
rect 793 321 797 325
rect 818 321 822 325
rect 954 321 958 325
rect 843 312 847 316
rect 1144 312 1148 316
rect 868 303 872 307
rect 1335 303 1339 307
rect 893 295 897 299
rect 1523 295 1527 299
rect 918 287 922 291
rect 1712 287 1716 291
rect 943 279 947 283
rect 1902 279 1906 283
rect 968 271 972 275
rect 2093 271 2097 275
rect 801 167 805 171
rect 826 158 830 162
rect 851 149 855 153
rect 876 141 880 145
rect 901 133 905 137
rect 926 125 930 129
rect 951 117 955 121
rect 976 109 980 113
rect 639 86 643 90
rect 698 2 702 6
<< metal2 >>
rect 639 372 643 603
rect 639 90 643 368
rect 698 6 702 687
rect 793 403 797 647
rect 801 526 805 647
rect 818 403 822 647
rect 826 535 830 647
rect 843 412 847 647
rect 851 544 855 647
rect 868 421 872 647
rect 876 552 880 647
rect 893 429 897 647
rect 901 560 905 647
rect 918 437 922 647
rect 926 568 930 647
rect 943 445 947 647
rect 951 576 955 647
rect 968 453 972 647
rect 976 584 980 647
rect 2044 494 2048 580
rect 2052 502 2056 572
rect 2060 510 2064 564
rect 2068 518 2072 556
rect 2076 526 2080 580
rect 2084 535 2088 572
rect 2092 544 2096 564
rect 2100 552 2104 556
rect 2108 518 2112 548
rect 2118 510 2122 540
rect 2127 502 2131 531
rect 2135 494 2139 522
rect 765 372 769 399
rect 765 325 769 368
rect 954 372 958 399
rect 793 325 797 331
rect 954 325 958 368
rect 793 46 797 321
rect 1144 372 1148 408
rect 801 46 805 167
rect 818 46 822 321
rect 1144 316 1148 368
rect 1335 372 1339 417
rect 826 46 830 158
rect 843 46 847 312
rect 1335 307 1339 368
rect 1523 372 1527 425
rect 851 46 855 149
rect 868 46 872 303
rect 1523 299 1527 368
rect 1712 372 1716 433
rect 876 46 880 141
rect 893 46 897 295
rect 1712 291 1716 368
rect 1902 372 1906 441
rect 901 46 905 133
rect 918 46 922 287
rect 1902 283 1906 368
rect 2093 372 2097 449
rect 926 46 930 125
rect 943 46 947 279
rect 2093 275 2097 368
rect 951 98 955 117
rect 968 46 972 271
rect 976 46 980 109
use BUFFER8  BUFFER8_1
timestamp 1746041965
transform 1 0 768 0 -1 90
box -4 -8 218 91
use BUFFER8  BUFFER8_0
timestamp 1746041965
transform 1 0 768 0 1 603
box -4 -8 218 91
<< labels >>
rlabel metal1 2265 169 2265 169 1 A0
rlabel metal1 2265 160 2265 160 1 A1
rlabel metal1 2265 151 2265 151 1 A2
rlabel metal1 2265 143 2265 143 1 A3
rlabel metal1 2265 135 2265 135 1 A4
rlabel metal1 2265 127 2265 127 1 A5
rlabel metal1 2265 119 2265 119 1 A6
rlabel metal1 2265 111 2265 111 1 A7
rlabel metal1 32 44 32 44 1 a_en
rlabel metal1 2262 524 2262 524 1 B7
rlabel metal1 2262 533 2262 533 1 B6
rlabel metal1 2262 542 2262 542 1 B5
rlabel metal1 2262 550 2262 550 1 B4
rlabel metal1 2262 558 2262 558 1 B3
rlabel metal1 2262 566 2262 566 1 B2
rlabel metal1 2262 574 2262 574 1 B1
rlabel metal1 2262 582 2262 582 1 B0
rlabel metal1 32 649 32 649 1 b_en
rlabel metal1 647 370 647 370 1 VSS
rlabel metal1 775 370 775 370 1 VSS
rlabel metal1 962 370 962 370 1 VSS
rlabel metal1 707 689 707 689 1 VDD
<< end >>
