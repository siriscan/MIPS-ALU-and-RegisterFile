magic
tech scmos
timestamp 1746041965
<< nwell >>
rect 0 260 14 264
rect 2187 260 2390 264
<< metal1 >>
rect 0 260 14 264
rect 2187 260 2390 264
rect 2066 224 2074 228
rect 2114 224 2122 228
rect 2070 220 2074 224
rect 2118 220 2122 224
rect 0 176 20 180
rect 2187 176 2272 180
rect 2276 176 2297 180
rect 2301 176 2322 180
rect 2326 176 2347 180
rect 2351 176 2372 180
rect 2376 176 2390 180
rect 2034 168 2062 172
rect 2082 160 2193 164
rect 2209 160 2388 164
rect 2018 152 2110 156
rect 2170 152 2222 156
rect 2234 152 2388 156
rect 2130 144 2247 148
rect 2259 144 2388 148
rect 2284 136 2388 140
rect 2309 128 2388 132
rect 2334 120 2388 124
rect 1920 112 2038 116
rect 2042 112 2086 116
rect 2090 112 2135 116
rect 2359 112 2388 116
rect 1000 104 1276 108
rect 2384 104 2388 108
rect 1016 96 1347 100
rect 9 88 13 92
rect 1000 88 1020 92
rect 9 80 13 84
rect 1008 80 1020 84
rect 9 72 13 76
rect 1016 72 1020 76
rect 9 64 13 68
rect 2 56 506 60
rect 2 48 514 52
rect 2 40 1012 44
rect 1351 40 2047 44
rect 2 32 1020 36
rect 6 24 10 28
rect 510 24 996 28
rect 1016 24 1020 28
rect 6 16 10 20
rect 518 16 1004 20
rect 6 8 10 12
rect 1280 8 2095 12
rect 6 0 10 4
rect 2 -8 1012 -4
rect 2 -16 1020 -12
rect 2 -24 1028 -20
rect 2 -32 1036 -28
rect 2 -40 890 -36
rect 902 -40 2143 -36
rect 894 -48 2174 -44
<< m2contact >>
rect 2062 210 2066 214
rect 2110 210 2114 214
rect 2047 206 2051 210
rect 2095 206 2099 210
rect 2143 209 2147 213
rect 2135 203 2139 207
rect 2038 196 2042 200
rect 2086 196 2090 200
rect 2272 192 2276 196
rect 2297 192 2301 196
rect 2322 192 2326 196
rect 2347 192 2351 196
rect 2372 192 2376 196
rect 2078 188 2082 192
rect 2126 188 2130 192
rect 2166 188 2170 192
rect 2272 176 2276 180
rect 2297 176 2301 180
rect 2322 176 2326 180
rect 2347 176 2351 180
rect 2372 176 2376 180
rect 2030 168 2034 172
rect 2062 168 2066 172
rect 2078 160 2082 164
rect 2193 160 2197 164
rect 2205 160 2209 164
rect 2014 152 2018 156
rect 2110 152 2114 156
rect 2166 152 2170 156
rect 2222 152 2226 156
rect 2230 152 2234 156
rect 2126 144 2130 148
rect 2247 144 2251 148
rect 2255 144 2259 148
rect 2280 136 2284 140
rect 2305 128 2309 132
rect 2330 120 2334 124
rect 1916 112 1920 116
rect 2038 112 2042 116
rect 2086 112 2090 116
rect 2135 112 2139 116
rect 2355 112 2359 116
rect 996 104 1000 108
rect 1276 104 1280 108
rect 2380 104 2384 108
rect 1012 96 1016 100
rect 1347 96 1351 100
rect 996 88 1000 92
rect 1004 80 1008 84
rect 1012 72 1016 76
rect 506 56 510 60
rect 514 48 518 52
rect 1012 40 1016 44
rect 1347 40 1351 44
rect 2047 40 2051 44
rect 1020 32 1024 36
rect 506 24 510 28
rect 996 24 1000 28
rect 1012 24 1016 28
rect 514 16 518 20
rect 1004 16 1008 20
rect 1020 16 1024 20
rect 1028 8 1032 12
rect 1276 8 1280 12
rect 2095 8 2099 12
rect 1012 -8 1016 -4
rect 1020 -16 1024 -12
rect 1028 -24 1032 -20
rect 1036 -32 1040 -28
rect 890 -40 894 -36
rect 898 -40 902 -36
rect 2143 -40 2147 -36
rect 890 -48 894 -44
rect 2174 -48 2178 -44
<< metal2 >>
rect 506 28 510 56
rect 514 20 518 48
rect 898 -36 902 116
rect 996 108 1000 116
rect 1012 100 1016 145
rect 2038 116 2042 196
rect 996 28 1000 88
rect 1004 20 1008 80
rect 1012 44 1016 72
rect 1020 36 1024 64
rect 1012 -4 1016 24
rect 1020 -12 1024 16
rect 1276 12 1280 104
rect 1347 44 1351 96
rect 2047 44 2051 206
rect 2062 172 2066 210
rect 2078 164 2082 188
rect 2086 116 2090 196
rect 2095 12 2099 206
rect 2110 156 2114 210
rect 2126 148 2130 188
rect 2135 116 2139 203
rect 1028 -20 1032 8
rect 1036 -28 1040 0
rect 2143 -36 2147 209
rect 2166 156 2170 188
rect 890 -44 894 -40
rect 2174 -44 2178 220
rect 2193 164 2197 216
rect 2205 164 2209 220
rect 2222 156 2226 220
rect 2230 156 2234 220
rect 2247 148 2251 220
rect 2255 148 2259 220
rect 2272 180 2276 192
rect 2280 140 2284 220
rect 2297 180 2301 192
rect 2305 132 2309 220
rect 2322 180 2326 192
rect 2330 124 2334 220
rect 2347 180 2351 192
rect 2355 116 2359 220
rect 2372 180 2376 192
rect 2380 108 2384 220
use AND2  AND2_0
timestamp 1740126148
transform 1 0 2132 0 1 176
box -5 0 45 92
use AOI21  AOI21_0
timestamp 1741232169
transform 1 0 2036 0 1 176
box -4 0 36 91
use AOI21  AOI21_1
timestamp 1741232169
transform 1 0 2084 0 1 176
box -4 0 36 91
use BUFFER8  BUFFER8_0
timestamp 1746041965
transform 1 0 2172 0 1 176
box -4 -8 218 91
use Comparator4  Comparator4_0
timestamp 1746041965
transform 1 0 0 0 1 136
box -4 -136 1022 132
use Comparator4  Comparator4_1
timestamp 1746041965
transform 1 0 1018 0 1 136
box -4 -136 1022 132
use INV  INV_0
timestamp 1741159900
transform 1 0 2068 0 1 176
box -4 0 20 91
use INV  INV_1
timestamp 1741159900
transform 1 0 2116 0 1 176
box -4 0 20 91
<< labels >>
rlabel metal1 10 90 10 90 1 A0
rlabel metal1 10 82 10 82 1 A1
rlabel metal1 10 74 10 74 1 A2
rlabel metal1 10 66 10 66 1 A3
rlabel metal1 10 58 10 58 1 A4
rlabel metal1 10 50 10 50 1 A5
rlabel metal1 10 42 10 42 1 A6
rlabel metal1 10 34 10 34 1 A7
rlabel metal1 7 26 7 26 1 B0
rlabel metal1 7 18 7 18 1 B1
rlabel metal1 7 10 7 10 1 B2
rlabel metal1 7 2 7 2 1 B3
rlabel metal1 7 -6 7 -6 1 B4
rlabel metal1 7 -14 7 -14 1 B5
rlabel metal1 7 -22 7 -22 1 B6
rlabel metal1 7 -30 7 -30 1 B7
rlabel metal1 5 -38 5 -38 1 enb
rlabel metal1 2386 162 2386 162 7 Y0
rlabel metal1 2386 154 2386 154 7 Y1
rlabel metal1 2386 146 2386 146 7 Y2
rlabel metal1 2386 138 2386 138 7 Y3
rlabel metal1 2386 130 2386 130 7 Y4
rlabel metal1 2386 122 2386 122 7 Y5
rlabel metal1 2386 114 2386 114 7 Y6
rlabel metal1 2386 106 2386 106 7 Y7
rlabel metal1 15 178 15 178 1 VSS
rlabel metal1 12 262 12 262 1 VDD
rlabel metal2 2168 173 2168 173 1 Equal
rlabel metal2 2080 169 2080 169 1 Less
rlabel metal2 2128 170 2128 170 1 Greater
<< end >>
