magic
tech scmos
timestamp 1746512792
<< nwell >>
rect -519 132 -516 136
rect -4 132 4 136
<< metal1 >>
rect -519 132 -516 136
rect -4 132 4 136
rect -519 48 -516 52
rect -4 48 4 52
rect -519 40 -514 44
rect -519 24 32 28
rect -531 0 -466 4
rect -454 0 23 4
rect -531 -8 -402 -4
rect -390 -8 212 -4
rect -531 -16 -338 -12
rect -326 -16 402 -12
rect -531 -24 -274 -20
rect -262 -24 593 -20
rect -531 -32 -210 -28
rect -198 -32 781 -28
rect -531 -40 -146 -36
rect -134 -40 970 -36
rect -531 -48 -82 -44
rect -70 -48 1160 -44
rect -531 -56 -18 -52
rect -6 -56 1351 -52
rect -531 -64 -491 -60
rect -487 -64 124 -60
rect 128 -64 1519 -60
rect -531 -72 -427 -68
rect -423 -72 313 -68
rect 317 -72 1519 -68
rect -531 -80 -363 -76
rect -359 -80 503 -76
rect 507 -80 1519 -76
rect -531 -88 -299 -84
rect -295 -88 694 -84
rect 698 -88 1519 -84
rect -531 -96 -235 -92
rect -231 -96 882 -92
rect 886 -96 1519 -92
rect -531 -104 -171 -100
rect -167 -104 1071 -100
rect 1075 -104 1519 -100
rect -531 -112 -107 -108
rect -103 -112 1261 -108
rect 1265 -112 1519 -108
rect -531 -120 -43 -116
rect -39 -120 1452 -116
rect 1456 -120 1519 -116
<< m2contact >>
rect 32 24 36 28
rect -466 0 -462 4
rect -458 0 -454 4
rect 23 0 27 4
rect -402 -8 -398 -4
rect -394 -8 -390 -4
rect 212 -8 216 -4
rect -338 -16 -334 -12
rect -330 -16 -326 -12
rect 402 -16 406 -12
rect -274 -24 -270 -20
rect -266 -24 -262 -20
rect 593 -24 597 -20
rect -210 -32 -206 -28
rect -202 -32 -198 -28
rect 781 -32 785 -28
rect -146 -40 -142 -36
rect -138 -40 -134 -36
rect 970 -40 974 -36
rect -82 -48 -78 -44
rect -74 -48 -70 -44
rect 1160 -48 1164 -44
rect -18 -56 -14 -52
rect -10 -56 -6 -52
rect 1351 -56 1355 -52
rect -491 -64 -487 -60
rect 124 -64 128 -60
rect -427 -72 -423 -68
rect 313 -72 317 -68
rect -363 -80 -359 -76
rect 503 -80 507 -76
rect -299 -88 -295 -84
rect 694 -88 698 -84
rect -235 -96 -231 -92
rect 882 -96 886 -92
rect -171 -104 -167 -100
rect 1071 -104 1075 -100
rect -107 -112 -103 -108
rect 1261 -112 1265 -108
rect -43 -120 -39 -116
rect 1452 -120 1456 -116
<< metal2 >>
rect -491 -60 -487 88
rect -466 4 -462 88
rect -458 4 -454 36
rect -427 -68 -423 88
rect -402 -4 -398 88
rect -394 -4 -390 32
rect -363 -76 -359 88
rect -338 -12 -334 88
rect -330 -12 -326 32
rect -299 -84 -295 88
rect -274 -20 -270 88
rect -266 -20 -262 32
rect -235 -92 -231 88
rect -210 -28 -206 88
rect -202 -28 -198 32
rect -171 -100 -167 88
rect -146 -36 -142 88
rect -138 -36 -134 32
rect -107 -108 -103 88
rect -82 -44 -78 88
rect -74 -44 -70 32
rect -43 -116 -39 88
rect -18 -52 -14 88
rect -10 -52 -6 32
rect 32 28 36 40
rect 124 -60 128 0
rect 212 -4 216 0
rect 313 -68 317 0
rect 402 -12 406 0
rect 503 -76 507 0
rect 593 -20 597 0
rect 694 -84 698 0
rect 781 -28 785 0
rect 882 -92 886 0
rect 970 -36 974 0
rect 1071 -100 1075 0
rect 1160 -44 1164 0
rect 1261 -108 1265 0
rect 1351 -52 1355 0
rect 1452 -116 1456 0
use 8bitMUX2to1  8bitMUX2to1_0
timestamp 1746042099
transform 1 0 -520 0 1 32
box 0 0 520 107
use reg8  reg8_0
timestamp 1745261002
transform 1 0 0 0 1 16
box 0 -16 1512 124
<< labels >>
rlabel metal1 -517 26 -517 26 3 clk
rlabel metal1 -517 42 -517 42 3 en
rlabel metal1 -529 2 -529 2 3 D0
rlabel metal1 -528 -6 -528 -6 3 D1
rlabel metal1 -528 -14 -528 -14 3 D2
rlabel metal1 -528 -22 -528 -22 3 D3
rlabel metal1 -528 -30 -528 -30 3 D4
rlabel metal1 -528 -38 -528 -38 3 D5
rlabel metal1 -528 -46 -528 -46 3 D6
rlabel metal1 -528 -54 -528 -54 3 D7
rlabel metal1 -517 50 -517 50 1 VSS
rlabel metal1 -518 134 -518 134 1 VDD
rlabel metal1 1517 -62 1517 -62 7 Q0
rlabel metal1 1517 -70 1517 -70 7 Q1
rlabel metal1 1516 -78 1516 -78 7 Q2
rlabel metal1 1516 -86 1516 -86 7 Q3
rlabel metal1 1516 -94 1516 -94 7 Q4
rlabel metal1 1516 -102 1516 -102 7 Q5
rlabel metal1 1517 -110 1517 -110 7 Q6
rlabel metal1 1516 -118 1516 -118 8 Q7
<< end >>
