magic
tech scmos
timestamp 1745340019
<< nwell >>
rect -6 44 125 96
<< ntransistor >>
rect 7 8 9 16
rect 15 8 17 16
rect 23 8 25 16
rect 39 8 41 12
rect 44 8 46 12
rect 62 8 64 12
rect 70 8 72 12
rect 78 8 80 12
rect 86 8 88 12
rect 102 8 104 12
rect 107 8 109 12
rect 112 8 114 12
<< ptransistor >>
rect 7 57 9 73
rect 15 57 17 73
rect 23 57 25 73
rect 39 69 41 73
rect 44 69 46 73
rect 62 69 64 73
rect 70 69 72 73
rect 78 69 80 73
rect 86 69 88 73
rect 102 69 104 73
rect 107 69 109 73
rect 112 69 114 73
<< ndiffusion >>
rect 6 8 7 16
rect 9 8 10 16
rect 14 8 15 16
rect 17 8 18 16
rect 22 8 23 16
rect 25 8 26 16
rect 38 8 39 12
rect 41 8 44 12
rect 46 8 47 12
rect 61 8 62 12
rect 64 8 65 12
rect 69 8 70 12
rect 72 8 73 12
rect 77 8 78 12
rect 80 8 81 12
rect 85 8 86 12
rect 88 8 89 12
rect 101 8 102 12
rect 104 8 107 12
rect 109 8 112 12
rect 114 8 115 12
<< pdiffusion >>
rect 6 57 7 73
rect 9 57 10 73
rect 14 57 15 73
rect 17 57 18 73
rect 22 57 23 73
rect 25 57 26 73
rect 38 69 39 73
rect 41 69 44 73
rect 46 69 47 73
rect 61 69 62 73
rect 64 69 65 73
rect 69 69 70 73
rect 72 69 73 73
rect 77 69 78 73
rect 80 69 81 73
rect 85 69 86 73
rect 88 69 89 73
rect 101 69 102 73
rect 104 69 107 73
rect 109 69 112 73
rect 114 69 115 73
<< ndcontact >>
rect 2 8 6 16
rect 10 8 14 16
rect 18 8 22 16
rect 26 8 30 16
rect 34 8 38 12
rect 47 8 51 12
rect 57 8 61 12
rect 65 8 69 12
rect 73 8 77 12
rect 81 8 85 12
rect 89 8 93 12
rect 97 8 101 12
rect 115 8 119 12
<< pdcontact >>
rect 2 57 6 73
rect 10 57 14 73
rect 18 57 22 73
rect 26 57 30 73
rect 34 69 38 73
rect 47 69 51 73
rect 57 69 61 73
rect 65 69 69 73
rect 73 69 77 73
rect 81 69 85 73
rect 89 69 93 73
rect 97 69 101 73
rect 115 69 119 73
<< psubstratepcontact >>
rect 10 0 14 4
rect 34 0 38 4
rect 57 0 61 4
rect 73 0 77 4
rect 97 0 101 4
<< nsubstratencontact >>
rect 10 84 14 88
rect 34 84 38 88
rect 57 84 61 88
rect 73 84 77 88
rect 97 84 101 88
<< polysilicon >>
rect 7 73 9 75
rect 15 73 17 75
rect 23 73 25 75
rect 39 73 41 75
rect 44 73 46 75
rect 62 73 64 75
rect 70 73 72 75
rect 78 73 80 75
rect 86 73 88 75
rect 102 73 104 75
rect 107 73 109 75
rect 112 73 114 75
rect 7 47 9 57
rect 8 43 9 47
rect 7 16 9 43
rect 15 40 17 57
rect 16 36 17 40
rect 14 26 16 36
rect 14 24 17 26
rect 15 16 17 24
rect 23 16 25 57
rect 39 47 41 69
rect 35 43 36 45
rect 40 43 41 47
rect 35 19 37 43
rect 35 17 41 19
rect 39 12 41 17
rect 44 12 46 69
rect 62 53 64 69
rect 63 49 64 53
rect 62 12 64 49
rect 70 45 72 69
rect 71 41 72 45
rect 70 12 72 41
rect 78 37 80 69
rect 79 33 80 37
rect 77 32 80 33
rect 77 22 79 32
rect 77 20 80 22
rect 78 12 80 20
rect 86 12 88 69
rect 102 40 104 69
rect 98 38 104 40
rect 98 16 100 38
rect 107 32 109 69
rect 103 21 105 31
rect 103 19 109 21
rect 98 14 104 16
rect 102 12 104 14
rect 107 12 109 19
rect 112 12 114 69
rect 7 6 9 8
rect 15 6 17 8
rect 23 6 25 8
rect 39 6 41 8
rect 44 6 46 8
rect 62 6 64 8
rect 70 6 72 8
rect 78 6 80 8
rect 86 6 88 8
rect 102 6 104 8
rect 107 6 109 8
rect 112 6 114 8
<< polycontact >>
rect 4 43 8 47
rect 12 36 16 40
rect 19 29 23 33
rect 36 43 40 47
rect 40 22 44 26
rect 59 49 63 53
rect 67 41 71 45
rect 75 33 79 37
rect 82 25 86 29
rect 98 43 102 47
rect 103 31 107 35
rect 108 24 112 28
<< metal1 >>
rect 0 84 10 88
rect 14 84 34 88
rect 38 84 57 88
rect 61 84 73 88
rect 77 84 97 88
rect 101 84 121 88
rect 10 73 14 84
rect 34 73 38 84
rect 57 73 61 84
rect 73 73 77 84
rect 97 73 101 84
rect 2 54 6 57
rect 18 54 22 57
rect 2 50 22 54
rect 2 19 22 23
rect 2 16 6 19
rect 18 16 22 19
rect 26 16 30 57
rect 47 12 51 69
rect 65 65 69 69
rect 81 65 85 69
rect 65 61 85 65
rect 89 63 93 69
rect 115 63 119 69
rect 89 59 119 63
rect 65 15 85 19
rect 65 12 69 15
rect 81 12 85 15
rect 89 12 93 59
rect 115 12 119 59
rect 10 4 14 8
rect 34 4 38 8
rect 57 4 61 8
rect 73 4 77 8
rect 97 4 101 8
rect 0 0 10 4
rect 14 0 34 4
rect 38 0 57 4
rect 61 0 73 4
rect 77 0 97 4
rect 101 0 121 4
rect -3 -8 51 -4
rect 55 -8 82 -4
rect 86 -8 116 -4
rect 8 -16 40 -12
rect 44 -16 59 -12
rect 63 -16 108 -12
rect 16 -24 32 -20
rect 36 -24 67 -20
rect 71 -24 99 -20
rect 23 -31 75 -27
rect 79 -31 90 -27
<< m2contact >>
rect 4 39 8 43
rect 12 40 16 44
rect 22 42 26 46
rect 19 33 23 37
rect 36 47 40 51
rect 40 26 44 30
rect 59 53 63 57
rect 67 45 71 49
rect 51 35 55 39
rect 75 37 79 41
rect 82 29 86 33
rect 98 47 102 51
rect 99 31 103 35
rect 108 20 112 24
rect 119 37 123 41
rect -7 -8 -3 -4
rect 51 -8 55 -4
rect 82 -8 86 -4
rect 4 -16 8 -12
rect 40 -16 44 -12
rect 59 -16 63 -12
rect 108 -16 112 -12
rect 12 -24 16 -20
rect 32 -24 36 -20
rect 67 -24 71 -20
rect 99 -24 103 -20
rect 19 -31 23 -27
rect 75 -31 79 -27
rect 90 -31 94 -27
<< metal2 >>
rect -7 50 26 54
rect -7 -4 -3 50
rect 4 43 8 47
rect 22 46 26 50
rect 4 -12 8 39
rect 12 -20 16 40
rect 19 -27 23 33
rect 32 -20 36 51
rect 40 -12 44 26
rect 51 -4 55 35
rect 59 -12 63 53
rect 67 -20 71 45
rect 90 47 98 51
rect 75 -27 79 37
rect 82 -4 86 29
rect 90 -27 94 47
rect 123 37 130 41
rect 103 31 107 35
rect 99 -20 103 31
rect 108 -12 112 20
<< labels >>
rlabel psubstratepcontact 12 2 12 2 1 VSS
rlabel metal1 83 -14 83 -14 1 A
rlabel metal1 52 -22 52 -22 1 B
rlabel metal1 52 -29 52 -29 1 C
rlabel metal2 128 39 128 39 1 Sb
rlabel nsubstratencontact 12 86 12 86 1 VDD
rlabel metal1 -1 -6 -1 -6 1 Cbout
<< end >>
