magic
tech scmos
timestamp 1740126148
<< nwell >>
rect -5 66 45 92
<< ntransistor >>
rect 7 8 9 16
rect 15 8 17 16
rect 31 8 33 12
<< ptransistor >>
rect 7 72 9 80
rect 15 72 17 80
rect 31 76 33 80
<< ndiffusion >>
rect 6 8 7 16
rect 9 8 15 16
rect 17 8 18 16
rect 30 8 31 12
rect 33 8 34 12
<< pdiffusion >>
rect 6 72 7 80
rect 9 72 10 80
rect 14 72 15 80
rect 17 72 18 80
rect 30 76 31 80
rect 33 76 34 80
<< ndcontact >>
rect 2 8 6 16
rect 18 8 22 16
rect 26 8 30 12
rect 34 8 38 12
<< pdcontact >>
rect 2 72 6 80
rect 10 72 14 80
rect 18 72 22 80
rect 26 76 30 80
rect 34 76 38 80
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 10 84 14 88
<< polysilicon >>
rect 7 80 9 82
rect 15 80 17 82
rect 31 80 33 82
rect 7 46 9 72
rect 4 44 9 46
rect 4 27 6 44
rect 7 16 9 27
rect 15 16 17 72
rect 31 12 33 76
rect 7 6 9 8
rect 15 6 17 8
rect 31 6 33 8
<< polycontact >>
rect 11 37 15 41
rect 3 23 7 27
rect 27 50 31 54
<< metal1 >>
rect 0 84 10 88
rect 14 84 40 88
rect 10 80 14 84
rect 26 80 30 84
rect 2 68 6 72
rect 18 68 22 72
rect 2 64 22 68
rect 18 54 22 64
rect 18 50 27 54
rect 18 16 22 50
rect 34 12 38 76
rect 2 4 6 8
rect 26 4 30 8
rect 0 0 2 4
rect 6 0 40 4
<< labels >>
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel nsubstratencontact 12 86 12 86 1 VDD
rlabel polycontact 5 25 5 25 1 B
rlabel polycontact 13 39 13 39 1 A
rlabel metal1 36 32 36 32 1 Y
<< end >>
