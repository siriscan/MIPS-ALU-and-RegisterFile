magic
tech scmos
timestamp 1746489366
<< metal1 >>
rect 20 120 24 124
rect 305 75 309 76
rect 15 36 19 40
rect 3400 36 3602 40
rect 3421 20 3600 24
rect -74 12 -33 16
rect 3446 12 3600 16
rect -38 4 117 8
rect 1142 4 1257 8
rect 2282 4 2397 8
rect 3471 4 3600 8
rect -74 -4 29 0
rect 33 -4 676 0
rect 1276 -4 2309 0
rect 2313 -4 2542 0
rect 2546 -4 3390 0
rect 3496 -4 3600 0
rect -74 -12 167 -8
rect 171 -12 814 -8
rect 1272 -12 1410 -8
rect 1414 -12 2334 -8
rect 2338 -12 2447 -8
rect 2451 -12 2680 -8
rect 2684 -12 3390 -8
rect 3521 -12 3600 -8
rect -74 -20 305 -16
rect 309 -20 952 -16
rect 1272 -20 1548 -16
rect 1552 -20 2472 -16
rect 2476 -20 2585 -16
rect 2589 -20 2818 -16
rect 2822 -20 3390 -16
rect 3546 -20 3600 -16
rect -74 -28 443 -24
rect 447 -28 1090 -24
rect 1272 -28 1686 -24
rect 1690 -28 2610 -24
rect 2614 -28 2723 -24
rect 2727 -28 2956 -24
rect 2960 -28 3390 -24
rect 3571 -28 3600 -24
rect -74 -36 54 -32
rect 58 -36 581 -32
rect 1272 -36 1824 -32
rect 1828 -36 2748 -32
rect 2752 -36 2861 -32
rect 2865 -36 3094 -32
rect 3098 -36 3390 -32
rect 3596 -36 3600 -32
rect -74 -44 192 -40
rect 196 -44 719 -40
rect 1272 -44 1962 -40
rect 1966 -44 2886 -40
rect 2890 -44 2999 -40
rect 3003 -44 3232 -40
rect 3236 -44 3390 -40
rect -74 -52 330 -48
rect 334 -52 857 -48
rect 1272 -52 2100 -48
rect 2104 -52 3024 -48
rect 3028 -52 3137 -48
rect 3141 -52 3370 -48
rect 3374 -52 3390 -48
rect -74 -60 -25 -56
rect -21 -60 468 -56
rect 472 -60 995 -56
rect 1272 -60 2238 -56
rect 2242 -60 3162 -56
rect 3166 -60 3275 -56
rect 3279 -60 3390 -56
rect 2 -68 606 -64
rect 610 -68 744 -64
rect 748 -68 882 -64
rect 886 -68 1020 -64
rect 1024 -68 2022 -64
rect 2026 -68 2160 -64
rect 2164 -68 3300 -64
rect -74 -76 -73 -72
rect -69 -76 1107 -72
rect 1111 -76 2247 -72
rect 2416 -80 3405 -76
rect -74 -84 2255 -80
rect 2259 -84 2286 -80
rect 2412 -88 2550 -84
rect 2554 -88 3434 -84
rect -74 -92 1115 -88
rect 1119 -92 1146 -88
rect 2412 -96 2688 -92
rect 2692 -96 3459 -92
rect -74 -100 -65 -96
rect -61 -100 6 -96
rect 136 -100 1169 -96
rect 1173 -100 1540 -96
rect 2412 -104 2826 -100
rect 2830 -104 3484 -100
rect 132 -108 270 -104
rect 274 -108 1307 -104
rect 1311 -108 1678 -104
rect 2412 -112 2964 -108
rect 2968 -112 3509 -108
rect 132 -116 408 -112
rect 412 -116 1194 -112
rect 1198 -116 1445 -112
rect 1449 -116 1816 -112
rect 2412 -120 3102 -116
rect 3106 -120 3534 -116
rect 132 -124 546 -120
rect 550 -124 1332 -120
rect 1336 -124 1583 -120
rect 1587 -124 1954 -120
rect 2412 -128 3240 -124
rect 3244 -128 3559 -124
rect 132 -132 684 -128
rect 688 -132 1470 -128
rect 1474 -132 1721 -128
rect 1725 -132 2092 -128
rect 2412 -136 3378 -132
rect 3382 -136 3584 -132
rect 132 -140 822 -136
rect 826 -140 1608 -136
rect 1612 -140 1859 -136
rect 1863 -140 2230 -136
rect 132 -148 960 -144
rect 964 -148 1746 -144
rect 1750 -148 1997 -144
rect 132 -156 1098 -152
rect 1102 -156 1884 -152
rect 1888 -156 2135 -152
rect -72 -164 3386 -160
<< m2contact >>
rect -65 69 -61 73
rect -25 69 -21 73
rect 1115 69 1119 73
rect 2255 69 2259 73
rect -73 55 -69 59
rect -33 55 -29 59
rect 1107 55 1111 59
rect 2247 55 2251 59
rect -42 48 -38 52
rect -2 48 2 52
rect 1138 48 1142 52
rect 2278 48 2282 52
rect 124 36 128 40
rect 262 36 266 40
rect 400 36 404 40
rect 538 36 542 40
rect 1264 36 1268 40
rect 1402 36 1406 40
rect 2404 36 2408 40
rect 3417 20 3421 24
rect -33 12 -29 16
rect 3442 12 3446 16
rect -42 4 -38 8
rect 1138 4 1142 8
rect 2278 4 2282 8
rect 3467 4 3471 8
rect 29 -4 33 0
rect 676 -4 680 0
rect 1272 -4 1276 0
rect 2309 -4 2313 0
rect 2542 -4 2546 0
rect 3492 -4 3496 0
rect 167 -12 171 -8
rect 814 -12 818 -8
rect 1410 -12 1414 -8
rect 2334 -12 2338 -8
rect 2447 -12 2451 -8
rect 2680 -12 2684 -8
rect 3517 -12 3521 -8
rect 305 -20 309 -16
rect 952 -20 956 -16
rect 1548 -20 1552 -16
rect 2472 -20 2476 -16
rect 2585 -20 2589 -16
rect 2818 -20 2822 -16
rect 3542 -20 3546 -16
rect 443 -28 447 -24
rect 1090 -28 1094 -24
rect 1686 -28 1690 -24
rect 2610 -28 2614 -24
rect 2723 -28 2727 -24
rect 2956 -28 2960 -24
rect 3567 -28 3571 -24
rect 54 -36 58 -32
rect 581 -36 585 -32
rect 1824 -36 1828 -32
rect 2748 -36 2752 -32
rect 2861 -36 2865 -32
rect 3094 -36 3098 -32
rect 3592 -36 3596 -32
rect 192 -44 196 -40
rect 719 -44 723 -40
rect 1962 -44 1966 -40
rect 2886 -44 2890 -40
rect 2999 -44 3003 -40
rect 3232 -44 3236 -40
rect 330 -52 334 -48
rect 857 -52 861 -48
rect 2100 -52 2104 -48
rect 3024 -52 3028 -48
rect 3137 -52 3141 -48
rect 3370 -52 3374 -48
rect -25 -60 -21 -56
rect 468 -60 472 -56
rect 995 -60 999 -56
rect 2238 -60 2242 -56
rect 3162 -60 3166 -56
rect 3275 -60 3279 -56
rect -2 -68 2 -64
rect 606 -68 610 -64
rect 744 -68 748 -64
rect 882 -68 886 -64
rect 1020 -68 1024 -64
rect 2022 -68 2026 -64
rect 2160 -68 2164 -64
rect 3300 -68 3304 -64
rect -73 -76 -69 -72
rect 1107 -76 1111 -72
rect 2247 -76 2251 -72
rect 2412 -80 2416 -76
rect 3405 -80 3409 -76
rect 2255 -84 2259 -80
rect 2286 -84 2290 -80
rect 2550 -88 2554 -84
rect 3434 -88 3438 -84
rect 1115 -92 1119 -88
rect 1146 -92 1150 -88
rect 2688 -96 2692 -92
rect 3459 -96 3463 -92
rect -65 -100 -61 -96
rect 6 -100 10 -96
rect 132 -100 136 -96
rect 1169 -100 1173 -96
rect 1540 -100 1544 -96
rect 2826 -104 2830 -100
rect 3484 -104 3488 -100
rect 270 -108 274 -104
rect 1307 -108 1311 -104
rect 1678 -108 1682 -104
rect 2964 -112 2968 -108
rect 3509 -112 3513 -108
rect 408 -116 412 -112
rect 1194 -116 1198 -112
rect 1445 -116 1449 -112
rect 1816 -116 1820 -112
rect 3102 -120 3106 -116
rect 3534 -120 3538 -116
rect 546 -124 550 -120
rect 1332 -124 1336 -120
rect 1583 -124 1587 -120
rect 1954 -124 1958 -120
rect 3240 -128 3244 -124
rect 3559 -128 3563 -124
rect 684 -132 688 -128
rect 1470 -132 1474 -128
rect 1721 -132 1725 -128
rect 2092 -132 2096 -128
rect 3378 -136 3382 -132
rect 3584 -136 3588 -132
rect 822 -140 826 -136
rect 1608 -140 1612 -136
rect 1859 -140 1863 -136
rect 2230 -140 2234 -136
rect 960 -148 964 -144
rect 1746 -148 1750 -144
rect 1997 -148 2001 -144
rect 1098 -156 1102 -152
rect 1884 -156 1888 -152
rect 2135 -156 2139 -152
rect 3386 -164 3390 -160
<< metal2 >>
rect -73 -72 -69 55
rect -65 -96 -61 69
rect -42 8 -38 48
rect -33 16 -29 55
rect -25 -56 -21 69
rect -2 -64 2 48
rect 6 -96 10 28
rect 29 0 33 76
rect 37 44 41 49
rect 54 -32 58 76
rect 107 44 111 49
rect 124 40 128 76
rect 132 -96 136 0
rect 167 -8 171 76
rect 175 44 179 49
rect 192 -40 196 76
rect 245 44 249 49
rect 262 40 266 76
rect 270 -104 274 0
rect 305 -16 309 76
rect 313 44 317 49
rect 330 -48 334 76
rect 383 44 387 52
rect 400 40 404 76
rect 408 -112 412 0
rect 443 -24 447 76
rect 451 44 455 49
rect 468 -56 472 76
rect 521 44 525 49
rect 538 40 542 76
rect 546 -120 550 0
rect 581 -32 585 76
rect 589 44 593 49
rect 606 -64 610 76
rect 659 44 663 49
rect 676 0 680 76
rect 684 -128 688 0
rect 719 -40 723 76
rect 727 44 731 49
rect 744 -64 748 76
rect 797 44 801 49
rect 814 -8 818 76
rect 822 -136 826 0
rect 857 -48 861 76
rect 865 44 869 49
rect 882 -64 886 76
rect 935 44 939 49
rect 952 -16 956 76
rect 960 -144 964 0
rect 995 -56 999 76
rect 1003 44 1007 49
rect 1020 -64 1024 76
rect 1073 44 1077 49
rect 1090 -24 1094 76
rect 1098 -152 1102 0
rect 1107 -72 1111 55
rect 1115 -88 1119 69
rect 1138 8 1142 48
rect 1146 -88 1150 28
rect 1169 -96 1173 76
rect 1177 44 1181 49
rect 1194 -112 1198 76
rect 1264 40 1268 76
rect 1272 0 1276 4
rect 1307 -104 1311 76
rect 1332 -120 1336 76
rect 1402 40 1406 76
rect 1410 -8 1414 4
rect 1445 -112 1449 76
rect 1470 -128 1474 76
rect 1540 -96 1544 80
rect 1548 -16 1552 4
rect 1583 -120 1587 76
rect 1608 -136 1612 76
rect 1678 -104 1682 76
rect 1686 -24 1690 4
rect 1721 -128 1725 76
rect 1746 -144 1750 76
rect 1816 -112 1820 76
rect 1824 -32 1828 4
rect 1859 -136 1863 76
rect 1884 -152 1888 76
rect 1954 -120 1958 76
rect 1962 -40 1966 4
rect 1997 -144 2001 76
rect 2022 -64 2026 76
rect 2092 -128 2096 76
rect 2100 -48 2104 4
rect 2135 -152 2139 76
rect 2160 -64 2164 76
rect 2230 -136 2234 76
rect 2238 -56 2242 4
rect 2247 -72 2251 55
rect 2255 -80 2259 69
rect 2278 8 2282 48
rect 2286 -80 2290 28
rect 2309 0 2313 76
rect 2334 -8 2338 76
rect 2404 40 2408 76
rect 2412 -76 2416 4
rect 2447 -8 2451 76
rect 2472 -16 2476 76
rect 2542 0 2546 76
rect 2550 -84 2554 4
rect 2585 -16 2589 76
rect 2610 -24 2614 76
rect 2680 -8 2684 76
rect 2688 -92 2692 4
rect 2723 -24 2727 76
rect 2748 -32 2752 76
rect 2818 -16 2822 76
rect 2826 -100 2830 4
rect 2861 -32 2865 76
rect 2886 -40 2890 76
rect 2956 -24 2960 76
rect 2964 -108 2968 4
rect 2999 -40 3003 76
rect 3024 -48 3028 76
rect 3094 -32 3098 76
rect 3102 -116 3106 4
rect 3137 -48 3141 76
rect 3162 -56 3166 76
rect 3232 -40 3236 76
rect 3240 -124 3244 4
rect 3275 -56 3279 76
rect 3300 -64 3304 76
rect 3370 -48 3374 76
rect 3378 -132 3382 4
rect 3386 -160 3390 80
rect 3405 -76 3409 76
rect 3417 24 3421 80
rect 3434 -84 3438 80
rect 3442 16 3446 80
rect 3459 -92 3463 80
rect 3467 8 3471 80
rect 3484 -100 3488 80
rect 3492 0 3496 80
rect 3509 -108 3513 80
rect 3517 -8 3521 80
rect 3534 -116 3538 80
rect 3542 -16 3546 80
rect 3559 -124 3563 80
rect 3567 -24 3571 80
rect 3584 -132 3588 80
rect 3592 -32 3596 80
use BUFFER8  BUFFER8_0
timestamp 1746041965
transform 1 0 3384 0 1 36
box -4 -8 218 91
use AND2  AND2_3
timestamp 1740126148
transform 1 0 2244 0 1 36
box -5 0 45 92
use AND2  AND2_2
timestamp 1740126148
transform 1 0 1104 0 1 36
box -5 0 45 92
use AND2  AND2_1
timestamp 1740126148
transform 1 0 -76 0 1 36
box -5 0 45 92
use AND2  AND2_0
timestamp 1740126148
transform 1 0 -36 0 1 36
box -5 0 45 92
use 8bitMUX3to1  8bitMUX3to1_0
timestamp 1746408420
transform 1 0 4 0 1 20
box -4 -20 1104 107
use 8bitMUX3to1  8bitMUX3to1_1
timestamp 1746408420
transform 1 0 1144 0 1 20
box -4 -20 1104 107
use 8bitMUX3to1  8bitMUX3to1_2
timestamp 1746408420
transform 1 0 2284 0 1 20
box -4 -20 1104 107
<< labels >>
rlabel metal1 17 38 17 38 1 VSS
rlabel metal1 22 122 22 122 5 VDD
rlabel metal1 -72 -2 -72 -2 1 A0
rlabel metal1 -72 -10 -72 -10 1 A1
rlabel metal1 -72 -18 -72 -18 1 A2
rlabel metal1 -72 -26 -72 -26 1 A3
rlabel metal1 -72 -34 -72 -34 1 A4
rlabel metal1 -72 -42 -72 -42 1 A5
rlabel metal1 -72 -50 -72 -50 1 A6
rlabel metal1 -72 -58 -72 -58 1 A7
rlabel metal1 -72 -82 -72 -82 1 B0
rlabel metal1 -72 -90 -72 -90 1 B1
rlabel metal1 -72 -98 -72 -98 1 B2
rlabel metal1 -67 14 -67 14 1 SIGN
rlabel metal1 -67 -74 -67 -74 1 RORL
rlabel metal1 -71 -162 -71 -162 1 ENb
rlabel metal1 138 -98 138 -98 1 first0
rlabel metal1 137 -106 137 -106 1 first1
rlabel metal1 137 -114 137 -114 1 first2
rlabel metal1 136 -122 136 -122 1 first3
rlabel metal1 136 -130 136 -130 1 first4
rlabel metal1 136 -138 136 -138 1 first5
rlabel metal1 136 -146 136 -146 1 first6
rlabel metal1 136 -154 136 -154 1 first7
rlabel metal1 1278 -2 1278 -2 1 second0
rlabel metal1 1278 -10 1278 -10 1 second1
rlabel metal1 1278 -18 1278 -18 1 second2
rlabel metal1 1278 -26 1278 -26 1 second3
rlabel metal1 1277 -34 1277 -34 1 second4
rlabel metal1 1277 -42 1277 -42 1 second5
rlabel metal1 1277 -50 1277 -50 1 second6
rlabel metal1 1276 -58 1276 -58 1 second7
rlabel metal1 3599 22 3599 22 7 Y0
rlabel metal1 3598 14 3598 14 7 Y1
rlabel metal1 3598 6 3598 6 7 Y2
rlabel metal1 3598 -2 3598 -2 7 Y3
rlabel metal1 3598 -10 3598 -10 7 Y4
rlabel metal1 3599 -18 3599 -18 7 Y5
rlabel metal1 3599 -26 3599 -26 7 Y6
rlabel metal1 3598 -34 3598 -34 7 Y7
<< end >>
