magic
tech scmos
timestamp 1746489366
<< nwell >>
rect 227 9074 231 9078
<< metal1 >>
rect 8 9153 7479 9157
rect 4 9145 12 9149
rect 16 9145 7487 9149
rect 4 9137 20 9141
rect 24 9137 7495 9141
rect 4 9129 28 9133
rect 32 9129 7503 9133
rect 4 9121 36 9125
rect 40 9121 7511 9125
rect 4 9113 44 9117
rect 48 9113 7519 9117
rect 4 9105 52 9109
rect 56 9105 7527 9109
rect 4 9097 60 9101
rect 64 9097 7535 9101
rect 227 9074 231 9078
rect -4 9034 0 9038
rect 1593 8931 1795 8935
rect 4 8821 8 8825
rect 4 8813 8 8817
rect 4 8805 8 8809
rect 4 8797 8 8801
rect 4 8789 8 8793
rect 4 8781 8 8785
rect 4 8773 8 8777
rect 4 8765 8 8769
rect 4 8180 16 8184
rect 4 8172 16 8176
rect 4 8164 16 8168
rect 4 8156 16 8160
rect 3351 8152 3352 8156
rect 3359 8152 3366 8156
rect 3359 8142 3366 8146
rect 3359 8133 3366 8137
rect 3359 8124 3366 8128
rect 3359 8116 3366 8120
rect 3359 8108 3366 8112
rect 3359 8100 3366 8104
rect 3359 8092 3366 8096
rect 0 8045 3379 8049
rect 0 8037 3371 8041
rect 0 8029 3363 8033
rect 3375 7880 3383 7884
rect 7531 7880 7543 7884
rect 3367 7872 3383 7876
rect 1569 7863 1574 7867
rect 3319 7841 3377 7845
rect 3311 7833 3377 7837
rect 3303 7825 3382 7829
rect 3295 7817 3382 7821
rect 3287 7809 3382 7813
rect 3279 7801 3382 7805
rect 3271 7793 3380 7797
rect 3263 7785 3378 7789
rect 3218 7777 3403 7781
rect 3210 7769 3403 7773
rect 5 7762 19 7766
rect 3202 7761 3403 7765
rect 5 7754 19 7758
rect 3194 7753 3403 7757
rect 5 7746 19 7750
rect 3186 7745 3403 7749
rect 3178 7737 3403 7741
rect 3170 7729 3403 7733
rect 3162 7721 3403 7725
rect 3360 7006 3363 7010
rect 3360 6996 3363 7000
rect 3360 6987 3363 6991
rect 3360 6978 3363 6982
rect 3360 6970 3363 6974
rect 3360 6962 3363 6966
rect 3360 6954 3363 6958
rect 3360 6946 3363 6950
rect 4 6736 22 6740
rect 4 6728 22 6732
rect 4 6720 22 6724
rect 0 6669 3377 6673
rect 0 6661 3377 6665
rect 3360 5832 3364 5836
rect 3360 5822 3364 5826
rect 3360 5813 3364 5817
rect 3360 5804 3364 5808
rect 3360 5796 3364 5800
rect 3360 5788 3364 5792
rect 3360 5780 3364 5784
rect 3360 5772 3364 5776
rect 3359 4660 3363 4664
rect 3359 4650 3363 4654
rect 3359 4641 3363 4645
rect 3359 4632 3363 4636
rect 3359 4624 3363 4628
rect 3359 4616 3363 4620
rect 3359 4608 3363 4612
rect 3359 4600 3363 4604
rect 3358 3501 3365 3505
rect 3358 3491 3365 3495
rect 3358 3482 3365 3486
rect 3358 3473 3365 3477
rect 3358 3465 3365 3469
rect 3358 3457 3365 3461
rect 3358 3449 3365 3453
rect 3358 3441 3365 3445
rect 3358 2345 3365 2349
rect 3358 2335 3365 2339
rect 3358 2326 3365 2330
rect 3358 2317 3365 2321
rect 3358 2309 3365 2313
rect 3358 2301 3365 2305
rect 3358 2293 3365 2297
rect 3358 2285 3365 2289
rect 3358 1187 3365 1191
rect 3358 1177 3365 1181
rect 3358 1168 3365 1172
rect 3358 1159 3365 1163
rect 3358 1151 3365 1155
rect 3358 1143 3365 1147
rect 3358 1135 3365 1139
rect 3358 1127 3365 1131
rect 3360 443 3365 447
rect 3358 433 3365 437
rect 3358 424 3365 428
rect 3358 415 3365 419
rect 3358 407 3365 411
rect 3358 399 3365 403
rect 3358 391 3365 395
rect 3358 383 3365 387
<< m2contact >>
rect 4 9153 8 9157
rect 7479 9153 7483 9157
rect 12 9145 16 9149
rect 7487 9145 7491 9149
rect 20 9137 24 9141
rect 7495 9137 7499 9141
rect 28 9129 32 9133
rect 7503 9129 7507 9133
rect 36 9121 40 9125
rect 7511 9121 7515 9125
rect 44 9113 48 9117
rect 7519 9113 7523 9117
rect 52 9105 56 9109
rect 7527 9105 7531 9109
rect 60 9097 64 9101
rect 7535 9097 7539 9101
rect 223 9074 227 9078
rect 4 8902 8 8906
rect 12 8894 16 8898
rect 20 8886 24 8890
rect 28 8878 32 8882
rect 36 8870 40 8874
rect 44 8862 48 8866
rect 52 8854 56 8858
rect 60 8845 64 8849
rect 3379 8045 3383 8049
rect 3371 8037 3375 8041
rect 3363 8029 3367 8033
rect 3379 7888 3383 7892
rect 3371 7880 3375 7884
rect 3363 7872 3367 7876
rect 3315 7841 3319 7845
rect 3307 7833 3311 7837
rect 3299 7825 3303 7829
rect 3291 7817 3295 7821
rect 3283 7809 3287 7813
rect 3275 7801 3279 7805
rect 3267 7793 3271 7797
rect 3259 7785 3263 7789
rect 3214 7777 3218 7781
rect 3206 7769 3210 7773
rect 3198 7761 3202 7765
rect 3190 7753 3194 7757
rect 3182 7745 3186 7749
rect 3174 7737 3178 7741
rect 3166 7729 3170 7733
rect 3158 7721 3162 7725
rect 3377 6688 3381 6692
rect 3377 6669 3381 6673
rect 3377 6661 3381 6665
rect 3377 6600 3381 6604
<< metal2 >>
rect 4 8906 8 9153
rect 12 8898 16 9145
rect 20 8890 24 9137
rect 28 8882 32 9129
rect 36 8874 40 9121
rect 44 8866 48 9113
rect 52 8858 56 9105
rect 60 8849 64 9097
rect 1608 8378 1612 8382
rect 3363 7876 3367 8029
rect 3371 7884 3375 8037
rect 3379 7892 3383 8045
rect 7479 7820 7483 9153
rect 7487 7820 7491 9145
rect 7495 7820 7499 9137
rect 7503 7820 7507 9129
rect 7511 7820 7515 9121
rect 7519 7820 7523 9113
rect 7527 7820 7531 9105
rect 7535 7820 7539 9097
rect 3158 7725 3162 7781
rect 3166 7733 3170 7781
rect 3166 7721 3170 7729
rect 3174 7741 3178 7781
rect 3174 7721 3178 7737
rect 3182 7749 3186 7781
rect 3182 7721 3186 7745
rect 3190 7757 3194 7781
rect 3190 7721 3194 7753
rect 3198 7765 3202 7781
rect 3198 7721 3202 7761
rect 3206 7773 3210 7781
rect 3206 7721 3210 7769
rect 3214 7721 3218 7777
rect 3377 6673 3381 6688
rect 3377 6604 3381 6661
rect 1448 197 1453 732
rect 3158 0 3162 1
rect 3166 0 3170 1
rect 3174 0 3178 1
rect 3182 0 3186 1
rect 3190 0 3194 1
rect 3198 0 3202 1
rect 3206 0 3210 1
rect 3214 0 3218 1
rect 3119 -4 3123 0
<< m3contact >>
rect 219 9074 223 9078
rect 1444 198 1448 202
<< metal3 >>
rect -1 9078 3393 9079
rect -1 9074 219 9078
rect 223 9074 3393 9078
rect -1 9073 3393 9074
rect 3387 7910 3393 9073
rect 3634 6419 3649 6425
rect 3634 203 3640 6419
rect -6 202 3640 203
rect -6 198 1444 202
rect 1448 198 3640 202
rect -6 197 3640 198
rect -6 196 1442 197
use ALU  ALU_0
timestamp 1746489366
transform 1 0 3794 0 1 6196
box -417 0 3745 1796
use REGISTER_FILE  REGISTER_FILE_0
timestamp 1746489366
transform 1 0 810 0 1 6666
box -810 -6666 2550 2428
<< labels >>
rlabel metal3 -3 200 -3 200 3 VSS
rlabel metal3 3 9076 3 9076 1 VDD
rlabel metal1 6 8823 6 8823 1 Imm0
rlabel metal1 6 8815 6 8815 1 Imm1
rlabel metal1 6 8807 6 8807 1 Imm2
rlabel metal1 6 8799 6 8799 1 Imm3
rlabel metal1 6 8791 6 8791 1 Imm4
rlabel metal1 6 8783 6 8783 1 Imm5
rlabel metal1 6 8775 6 8775 1 Imm6
rlabel metal1 6 8767 6 8767 1 Imm7
rlabel metal1 7468 9155 7468 9155 7 Y0
rlabel metal1 7467 9147 7467 9147 7 Y1
rlabel metal1 7467 9139 7467 9139 7 Y2
rlabel metal1 7466 9131 7466 9131 7 Y3
rlabel metal1 7467 9123 7467 9123 7 Y4
rlabel metal1 7467 9115 7467 9115 7 Y5
rlabel metal1 7467 9107 7467 9107 7 Y6
rlabel metal1 7467 9099 7467 9099 1 Y7
rlabel metal1 7541 7882 7541 7882 7 Overflow
rlabel metal1 9 8182 9 8182 1 Write_Address0
rlabel metal1 9 8174 9 8174 1 Write_Address1
rlabel metal1 9 8166 9 8166 1 Write_Address2
rlabel metal1 9 8158 9 8158 1 Write_Address3
rlabel metal1 10 7764 10 7764 1 B_Read_Address0
rlabel metal1 8 7756 8 7756 1 B_Read_Address1
rlabel metal1 10 7748 10 7748 1 B_Read_Address2
rlabel metal1 11 6738 11 6738 1 A_Read_Address0
rlabel metal1 10 6730 10 6730 1 A_Read_Address1
rlabel metal1 10 6722 10 6722 1 A_Read_Address2
rlabel metal1 0 8047 0 8047 3 func0
rlabel metal1 0 8039 0 8039 3 func1
rlabel metal1 0 8031 0 8031 3 func2
rlabel metal1 3 6663 3 6663 1 RorL
rlabel metal1 2 6671 2 6671 1 LorA
rlabel metal1 3364 8154 3364 8154 1 reg_zero0
rlabel metal1 3364 8144 3364 8144 1 reg_zero1
rlabel metal1 3364 8135 3364 8135 1 reg_zero2
rlabel metal1 3363 8126 3363 8126 1 reg_zero3
rlabel metal1 3361 8118 3361 8118 1 reg_zero4
rlabel metal1 3361 8110 3361 8110 1 reg_zero5
rlabel metal1 3361 8102 3361 8102 1 reg_zero6
rlabel metal1 3362 8094 3362 8094 1 reg_zero7
rlabel metal1 -2 9036 -2 9036 3 imm_en
rlabel metal1 3361 7008 3361 7008 1 reg_one0
rlabel metal1 3361 6998 3361 6998 1 reg_one1
rlabel metal1 3361 6989 3361 6989 1 reg_one2
rlabel metal1 3361 6980 3361 6980 1 reg_one3
rlabel metal1 3361 6972 3361 6972 1 reg_one4
rlabel metal1 3361 6964 3361 6964 1 reg_one5
rlabel metal1 3361 6956 3361 6956 1 reg_one6
rlabel metal1 3361 6948 3361 6948 1 reg_one7
rlabel metal1 3361 5834 3361 5834 1 reg_two0
rlabel metal1 3361 5824 3361 5824 1 reg_two1
rlabel metal1 3361 5815 3361 5815 1 reg_two2
rlabel metal1 3361 5806 3361 5806 1 reg_two3
rlabel metal1 3361 5798 3361 5798 1 reg_two4
rlabel metal1 3361 5790 3361 5790 1 reg_two5
rlabel metal1 3361 5782 3361 5782 1 reg_two6
rlabel metal1 3361 5774 3361 5774 1 reg_two7
rlabel metal1 3361 4662 3361 4662 1 reg_three0
rlabel metal1 3361 4652 3361 4652 1 reg_three1
rlabel metal1 3362 4643 3362 4643 1 reg_three2
rlabel metal1 3362 4634 3362 4634 1 reg_three3
rlabel metal1 3362 4626 3362 4626 1 reg_three4
rlabel metal1 3362 4618 3362 4618 1 reg_three5
rlabel metal1 3362 4610 3362 4610 1 reg_three6
rlabel metal1 3362 4602 3362 4602 1 reg_three7
rlabel metal1 3361 3503 3361 3503 1 reg_four0
rlabel metal1 3362 3493 3362 3493 1 reg_four1
rlabel metal1 3362 3484 3362 3484 1 reg_four2
rlabel metal1 3362 3475 3362 3475 1 reg_four3
rlabel metal1 3362 3467 3362 3467 1 reg_four4
rlabel metal1 3362 3459 3362 3459 1 reg_four5
rlabel metal1 3362 3451 3362 3451 1 reg_four6
rlabel metal1 3362 3443 3362 3443 1 reg_four7
rlabel metal1 3362 2347 3362 2347 1 reg_five0
rlabel metal1 3362 2337 3362 2337 1 reg_five1
rlabel metal1 3362 2328 3362 2328 1 reg_five2
rlabel metal1 3362 2319 3362 2319 1 reg_five3
rlabel metal1 3362 2311 3362 2311 1 reg_five4
rlabel metal1 3362 2303 3362 2303 1 reg_five5
rlabel metal1 3362 2295 3362 2295 1 reg_five6
rlabel metal1 3362 2287 3362 2287 1 reg_five7
rlabel metal1 3362 1189 3362 1189 1 reg_six0
rlabel metal1 3362 1179 3362 1179 1 reg_six1
rlabel metal1 3362 1170 3362 1170 1 reg_six2
rlabel metal1 3362 1161 3362 1161 1 reg_six3
rlabel metal1 3361 1153 3361 1153 1 reg_six4
rlabel metal1 3361 1145 3361 1145 1 reg_six5
rlabel metal1 3361 1137 3361 1137 1 reg_six6
rlabel metal1 3362 1129 3362 1129 1 reg_six7
rlabel metal2 3121 -2 3121 -2 1 clk
rlabel metal2 1610 8380 1610 8380 1 check
rlabel metal1 3325 7843 3325 7843 3 A0
rlabel metal1 3325 7835 3325 7835 3 A1
rlabel metal1 3325 7827 3325 7827 3 A2
rlabel metal1 3325 7819 3325 7819 3 A3
rlabel metal1 3325 7811 3325 7811 3 A4
rlabel metal1 3325 7803 3325 7803 3 A5
rlabel metal1 3325 7795 3325 7795 3 A6
rlabel metal1 3325 7787 3325 7787 3 A7
rlabel metal1 3325 7779 3325 7779 3 B0
rlabel metal1 3325 7771 3325 7771 3 B1
rlabel metal1 3325 7763 3325 7763 3 B2
rlabel metal1 3325 7755 3325 7755 3 B3
rlabel metal1 3325 7747 3325 7747 3 B4
rlabel metal1 3325 7739 3325 7739 3 B5
rlabel metal1 3325 7731 3325 7731 3 B6
rlabel metal1 3325 7723 3325 7723 3 B7
rlabel metal1 1571 7865 1571 7865 1 D0
rlabel metal1 3361 445 3361 445 1 reg_seven
<< end >>
