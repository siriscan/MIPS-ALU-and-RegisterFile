magic
tech scmos
timestamp 1746041965
<< nwell >>
rect 2135 121 2337 125
<< metal1 >>
rect 10 121 14 125
rect 2135 121 2337 125
rect 2006 77 2010 81
rect 453 69 457 73
rect 22 57 26 67
rect 245 57 249 61
rect 273 57 277 67
rect 364 61 368 65
rect 321 59 325 60
rect 524 57 528 67
rect 321 53 325 57
rect 775 57 779 67
rect 1026 57 1030 67
rect 1277 57 1281 67
rect 1528 57 1532 67
rect 1779 57 1783 67
rect 2026 57 2030 67
rect 10 37 14 41
rect 2135 37 2337 41
rect 203 29 237 33
rect 453 29 488 33
rect 705 29 739 33
rect 956 29 990 33
rect 1207 29 1241 33
rect 1458 29 1492 33
rect 1709 29 1743 33
rect 1960 29 1994 33
rect 2078 29 2105 33
rect 2117 21 2335 25
rect 2156 13 2335 17
rect 10 6 106 10
rect 249 6 357 10
rect 500 6 608 10
rect 751 6 859 10
rect 1002 6 1110 10
rect 1253 6 1361 10
rect 1504 6 1613 10
rect 1755 6 1863 10
rect 2181 5 2335 9
rect 181 -2 257 2
rect 261 -2 508 2
rect 512 -2 759 2
rect 763 -2 1010 2
rect 1014 -2 1261 2
rect 1265 -2 1512 2
rect 1516 -2 1763 2
rect 1767 -2 2026 2
rect 2206 -3 2335 1
rect 6 -10 2082 -6
rect 2231 -11 2335 -7
rect 6 -18 91 -14
rect 233 -18 2140 -14
rect 2256 -19 2335 -15
rect 6 -26 342 -22
rect 484 -26 2169 -22
rect 2281 -27 2335 -23
rect 6 -34 593 -30
rect 735 -34 2194 -30
rect 2306 -35 2335 -31
rect 6 -42 844 -38
rect 986 -42 2219 -38
rect 2331 -43 2335 -39
rect 6 -50 1095 -46
rect 1237 -50 2244 -46
rect 6 -58 1346 -54
rect 1488 -58 2269 -54
rect 6 -66 1597 -62
rect 1739 -66 2294 -62
rect 6 -74 1848 -70
rect 1990 -74 2319 -70
rect 6 -82 22 -78
rect 6 -90 273 -86
rect 6 -98 524 -94
rect 6 -106 775 -102
rect 6 -114 1026 -110
rect 6 -122 1277 -118
rect 6 -130 1528 -126
rect 6 -138 1779 -134
<< m2contact >>
rect 237 73 241 77
rect 488 73 492 77
rect 739 73 743 77
rect 990 73 994 77
rect 1241 73 1245 77
rect 1492 73 1496 77
rect 1743 73 1747 77
rect 1994 73 1998 77
rect 22 53 26 57
rect 273 53 277 57
rect 524 53 528 57
rect 775 53 779 57
rect 1026 53 1030 57
rect 1277 53 1281 57
rect 1528 53 1532 57
rect 1779 53 1783 57
rect 2026 53 2030 57
rect 229 49 233 53
rect 245 49 249 53
rect 480 49 484 53
rect 496 49 500 53
rect 731 49 735 53
rect 747 49 751 53
rect 982 49 986 53
rect 998 49 1002 53
rect 1233 49 1237 53
rect 1249 49 1253 53
rect 1484 49 1488 53
rect 1500 49 1504 53
rect 1735 49 1739 53
rect 1751 49 1755 53
rect 1986 49 1990 53
rect 2074 49 2078 53
rect 237 29 241 33
rect 488 29 492 33
rect 739 29 743 33
rect 990 29 994 33
rect 1241 29 1245 33
rect 1492 29 1496 33
rect 1743 29 1747 33
rect 1994 29 1998 33
rect 2074 29 2078 33
rect 2105 29 2109 33
rect 2113 21 2117 25
rect 2152 13 2156 17
rect 6 6 10 10
rect 245 6 249 10
rect 496 6 500 10
rect 747 6 751 10
rect 998 6 1002 10
rect 1249 6 1253 10
rect 1500 6 1504 10
rect 1751 6 1755 10
rect 2177 5 2181 9
rect 177 -2 181 2
rect 257 -2 261 2
rect 508 -2 512 2
rect 759 -2 763 2
rect 1010 -2 1014 2
rect 1261 -2 1265 2
rect 1512 -2 1516 2
rect 1763 -2 1767 2
rect 2026 -2 2030 2
rect 2202 -3 2206 1
rect 2082 -10 2086 -6
rect 2227 -11 2231 -7
rect 91 -18 95 -14
rect 229 -18 233 -14
rect 2140 -18 2144 -14
rect 2252 -19 2256 -15
rect 342 -26 346 -22
rect 480 -26 484 -22
rect 2169 -26 2173 -22
rect 2277 -27 2281 -23
rect 593 -34 597 -30
rect 731 -34 735 -30
rect 2194 -34 2198 -30
rect 2302 -35 2306 -31
rect 844 -42 848 -38
rect 982 -42 986 -38
rect 2219 -42 2223 -38
rect 2327 -43 2331 -39
rect 1095 -50 1099 -46
rect 1233 -50 1237 -46
rect 2244 -50 2248 -46
rect 1346 -58 1350 -54
rect 1484 -58 1488 -54
rect 2269 -58 2273 -54
rect 1597 -66 1601 -62
rect 1735 -66 1739 -62
rect 2294 -66 2298 -62
rect 1848 -74 1852 -70
rect 1986 -74 1990 -70
rect 2319 -74 2323 -70
rect 22 -82 26 -78
rect 273 -90 277 -86
rect 524 -98 528 -94
rect 775 -106 779 -102
rect 1026 -114 1030 -110
rect 1277 -122 1281 -118
rect 1528 -130 1532 -126
rect 1779 -138 1783 -134
<< metal2 >>
rect 2086 81 2121 85
rect 6 10 10 60
rect 22 -78 26 53
rect 91 -14 95 21
rect 177 2 181 6
rect 229 -14 233 49
rect 237 33 241 73
rect 245 10 249 49
rect 257 2 261 60
rect 273 -86 277 53
rect 342 -22 346 29
rect 480 -22 484 49
rect 488 33 492 73
rect 496 10 500 49
rect 508 2 512 60
rect 524 -94 528 53
rect 593 -30 597 21
rect 731 -30 735 49
rect 739 33 743 73
rect 747 10 751 49
rect 759 2 763 60
rect 775 -102 779 53
rect 844 -38 848 21
rect 982 -38 986 49
rect 990 33 994 73
rect 998 10 1002 49
rect 1010 2 1014 60
rect 1026 -110 1030 53
rect 1095 -46 1099 21
rect 1233 -46 1237 49
rect 1241 33 1245 73
rect 1249 10 1253 49
rect 1261 2 1265 60
rect 1277 -118 1281 53
rect 1346 -54 1350 25
rect 1484 -54 1488 49
rect 1492 33 1496 73
rect 1500 10 1504 49
rect 1512 2 1516 60
rect 1528 -126 1532 53
rect 1597 -62 1601 25
rect 1735 -62 1739 49
rect 1743 33 1747 73
rect 1751 10 1755 49
rect 1763 2 1767 60
rect 1779 -134 1783 53
rect 1848 -70 1852 25
rect 1986 -70 1990 49
rect 1994 33 1998 73
rect 2026 2 2030 53
rect 2074 33 2078 49
rect 2082 -6 2086 81
rect 2105 33 2109 73
rect 2113 25 2117 73
rect 2140 -14 2144 77
rect 2152 17 2156 81
rect 2169 -22 2173 81
rect 2177 9 2181 81
rect 2194 -30 2198 81
rect 2202 1 2206 81
rect 2219 -38 2223 81
rect 2227 -7 2231 81
rect 2244 -46 2248 81
rect 2252 -15 2256 81
rect 2269 -54 2273 81
rect 2277 -23 2281 81
rect 2294 -62 2298 81
rect 2302 -31 2306 81
rect 2319 -70 2323 81
rect 2327 -39 2331 81
use 1bitAddSub  1bitAddSub_0
timestamp 1746041965
transform 1 0 80 0 1 0
box -80 6 159 133
use INV  INV_0
timestamp 1741159900
transform 1 0 235 0 1 37
box -4 0 20 91
use 1bitAddSub  1bitAddSub_1
timestamp 1746041965
transform 1 0 331 0 1 0
box -80 6 159 133
use 1bitAddSub  1bitAddSub_2
timestamp 1746041965
transform 1 0 582 0 1 0
box -80 6 159 133
use INV  INV_1
timestamp 1741159900
transform 1 0 486 0 1 37
box -4 0 20 91
use 1bitAddSub  1bitAddSub_3
timestamp 1746041965
transform 1 0 833 0 1 0
box -80 6 159 133
use INV  INV_2
timestamp 1741159900
transform 1 0 737 0 1 37
box -4 0 20 91
use 1bitAddSub  1bitAddSub_4
timestamp 1746041965
transform 1 0 1084 0 1 0
box -80 6 159 133
use INV  INV_3
timestamp 1741159900
transform 1 0 988 0 1 37
box -4 0 20 91
use 1bitAddSub  1bitAddSub_5
timestamp 1746041965
transform 1 0 1335 0 1 0
box -80 6 159 133
use INV  INV_4
timestamp 1741159900
transform 1 0 1239 0 1 37
box -4 0 20 91
use 1bitAddSub  1bitAddSub_6
timestamp 1746041965
transform 1 0 1586 0 1 0
box -80 6 159 133
use INV  INV_5
timestamp 1741159900
transform 1 0 1490 0 1 37
box -4 0 20 91
use 1bitAddSub  1bitAddSub_7
timestamp 1746041965
transform 1 0 1837 0 1 0
box -80 6 159 133
use INV  INV_6
timestamp 1741159900
transform 1 0 1741 0 1 37
box -4 0 20 91
use BUFFER8  BUFFER8_0
timestamp 1746041965
transform 1 0 2119 0 1 37
box -4 -8 218 91
use BUFFER  BUFFER_0
timestamp 1746041965
transform 1 0 2080 0 1 37
box -4 0 43 91
use INV  INV_7
timestamp 1741159900
transform 1 0 1992 0 1 37
box -4 0 20 91
use XOR2  XOR2_0
timestamp 1746041965
transform 1 0 2040 0 1 37
box -36 0 44 94
<< labels >>
rlabel metal1 12 8 12 8 1 K
rlabel metal1 8 -8 8 -8 1 enb
rlabel metal1 12 123 12 123 1 VDD
rlabel metal1 12 39 12 39 1 VSS
rlabel metal1 8 -80 8 -80 1 B0
rlabel metal1 8 -88 8 -88 1 B1
rlabel metal1 8 -96 8 -96 1 B2
rlabel metal1 8 -104 8 -104 1 B3
rlabel metal1 8 -112 8 -112 1 B4
rlabel metal1 8 -120 8 -120 1 B5
rlabel metal1 8 -128 8 -128 1 B6
rlabel metal1 8 -136 8 -136 1 B7
rlabel metal1 8 -16 8 -16 1 A0
rlabel metal1 8 -24 8 -24 1 A1
rlabel metal1 8 -32 8 -32 1 A2
rlabel metal1 8 -40 8 -40 1 A3
rlabel metal1 8 -48 8 -48 1 A4
rlabel metal1 8 -56 8 -56 1 A5
rlabel metal1 8 -64 8 -64 1 A6
rlabel metal1 8 -72 8 -72 1 A7
rlabel metal1 2333 23 2333 23 1 Overflow
rlabel metal1 2333 15 2333 15 1 D0
rlabel metal1 2333 7 2333 7 1 D1
rlabel metal1 2333 -1 2333 -1 1 D2
rlabel metal1 2333 -9 2333 -9 1 D3
rlabel metal1 2333 -17 2333 -17 1 D4
rlabel metal1 2333 -25 2333 -25 1 D5
rlabel metal1 2333 -33 2333 -33 1 D6
rlabel metal1 2333 -41 2333 -41 1 D7
<< end >>
