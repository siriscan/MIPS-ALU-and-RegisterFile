magic
tech scmos
timestamp 1746489366
<< nwell >>
rect -583 2427 715 2428
rect -583 2389 716 2427
rect 684 2278 716 2389
rect -245 1652 -192 1677
rect -209 1624 -192 1652
rect -209 1606 117 1624
rect -281 1312 715 1338
rect -281 1236 -257 1312
rect 684 1134 709 1147
rect 96 254 123 316
rect -300 226 123 254
rect 684 -40 712 3
rect 684 -1216 715 -1172
rect 684 -2371 710 -2346
rect 684 -3527 711 -3505
rect 684 -4685 709 -4661
rect 684 -5819 710 -5818
rect 684 -5859 712 -5819
<< metal1 >>
rect -67 2408 697 2412
rect -810 2368 -577 2372
rect -67 2324 638 2328
rect -517 2301 -19 2305
rect -453 2293 -27 2297
rect -389 2285 -35 2289
rect -325 2277 -43 2281
rect -261 2269 -51 2273
rect -197 2261 -59 2265
rect -133 2253 -66 2257
rect -810 2236 -554 2240
rect -810 2228 -490 2232
rect -5 2225 32 2229
rect -810 2220 -426 2224
rect -810 2212 -362 2216
rect -810 2204 -298 2208
rect -810 2196 -234 2200
rect -810 2188 -170 2192
rect -810 2179 -106 2183
rect -810 2155 -529 2159
rect 2263 2158 2404 2162
rect -810 2147 -465 2151
rect 2263 2150 2396 2154
rect -810 2139 -401 2143
rect 2263 2142 2388 2146
rect -810 2131 -337 2135
rect 2263 2134 2380 2138
rect -810 2123 -273 2127
rect 2263 2126 2372 2130
rect -810 2115 -209 2119
rect 2263 2118 2364 2122
rect -810 2107 -145 2111
rect 2263 2109 2356 2113
rect -810 2099 -81 2103
rect 2254 2100 2348 2104
rect -169 1911 -9 1915
rect -15 1732 0 1736
rect -23 1723 0 1727
rect -31 1715 0 1719
rect -39 1707 0 1711
rect -47 1699 0 1703
rect -55 1691 0 1695
rect -62 1683 0 1687
rect -69 1675 0 1679
rect -249 1670 -204 1674
rect -200 1617 112 1621
rect -249 1586 13 1590
rect -810 1514 -751 1518
rect -810 1506 -735 1510
rect -810 1498 -719 1502
rect -810 1490 -767 1494
rect 2138 1486 2550 1490
rect 2138 1476 2550 1480
rect 2138 1467 2550 1471
rect 2138 1458 2550 1462
rect -363 1453 30 1457
rect 2138 1450 2550 1454
rect -347 1445 -99 1449
rect 2138 1442 2550 1446
rect -331 1437 -106 1441
rect 2138 1434 2550 1438
rect -315 1429 -114 1433
rect 2138 1426 2550 1430
rect -299 1421 -122 1425
rect -283 1413 -130 1417
rect -267 1405 -138 1409
rect 2188 1387 2309 1391
rect -267 1325 697 1329
rect 2266 1322 2505 1326
rect 2266 1313 2497 1317
rect 2266 1304 2489 1308
rect 2266 1296 2481 1300
rect 2266 1288 2473 1292
rect 2266 1280 2465 1284
rect 2266 1272 2457 1276
rect 2266 1264 2449 1268
rect -276 1252 -271 1256
rect 17 1241 648 1245
rect -250 1197 33 1201
rect -672 1168 -666 1172
rect -276 1168 13 1172
rect -672 1156 -666 1160
rect -810 1096 -650 1100
rect -810 1088 -634 1092
rect -565 1087 -173 1091
rect -810 1080 -618 1084
rect -524 1079 33 1083
rect -483 1071 -189 1075
rect -442 1063 -197 1067
rect -401 1055 -205 1059
rect -360 1047 -213 1051
rect -319 1039 -220 1043
rect -278 1031 -227 1035
rect 2263 1012 2404 1016
rect 2263 1004 2396 1008
rect 2263 996 2388 1000
rect 2263 988 2380 992
rect 2263 980 2372 984
rect 2263 972 2364 976
rect 2263 963 2356 967
rect 2263 954 2348 958
rect -15 586 0 590
rect -23 577 0 581
rect -31 569 0 573
rect -39 561 0 565
rect -47 553 0 557
rect -55 545 0 549
rect -62 537 0 541
rect -69 529 0 533
rect 2264 340 2550 344
rect 2264 330 2550 334
rect 2264 321 2550 325
rect 2264 312 2550 316
rect -95 307 32 311
rect 2264 304 2550 308
rect 2264 296 2550 300
rect 2264 288 2550 292
rect 2264 280 2550 284
rect -302 242 112 246
rect 2264 241 2309 245
rect 2266 176 2505 180
rect 2266 167 2497 171
rect -698 158 -694 162
rect -302 158 638 162
rect 2266 158 2489 162
rect 2266 150 2481 154
rect -698 146 -692 150
rect 2266 142 2473 146
rect 2266 134 2465 138
rect 2266 126 2457 130
rect 2266 118 2449 122
rect -810 70 -676 74
rect -810 62 -660 66
rect -591 59 -254 63
rect -810 54 -644 58
rect -550 51 29 55
rect -509 43 -270 47
rect -468 35 -278 39
rect -427 27 -286 31
rect -386 19 -294 23
rect -345 11 -301 15
rect -185 -95 33 -91
rect 2263 -162 2404 -158
rect 2263 -170 2396 -166
rect 2263 -178 2388 -174
rect 2263 -186 2380 -182
rect 2263 -194 2372 -190
rect 2263 -202 2364 -198
rect 2263 -211 2356 -207
rect 2263 -220 2348 -216
rect -15 -588 0 -584
rect -23 -597 0 -593
rect -31 -605 0 -601
rect -39 -613 0 -609
rect -47 -621 0 -617
rect -55 -629 0 -625
rect -62 -637 0 -633
rect -69 -645 0 -641
rect 2257 -834 2550 -830
rect 2257 -844 2550 -840
rect 2257 -853 2550 -849
rect 2257 -862 2550 -858
rect -102 -867 30 -863
rect 2257 -870 2550 -866
rect 2257 -878 2550 -874
rect 2257 -886 2550 -882
rect 2257 -894 2550 -890
rect 2264 -933 2309 -929
rect 2266 -998 2505 -994
rect 2266 -1007 2497 -1003
rect 2266 -1016 2489 -1012
rect 2266 -1024 2481 -1020
rect 2266 -1032 2473 -1028
rect 2266 -1040 2465 -1036
rect 2266 -1048 2457 -1044
rect 2266 -1056 2449 -1052
rect -266 -1123 32 -1119
rect -193 -1267 33 -1263
rect 2263 -1334 2404 -1330
rect 2263 -1342 2396 -1338
rect 2263 -1350 2388 -1346
rect 2263 -1358 2380 -1354
rect 2263 -1366 2372 -1362
rect 2263 -1374 2364 -1370
rect 2263 -1383 2356 -1379
rect 2263 -1392 2348 -1388
rect -15 -1760 2 -1756
rect -23 -1769 2 -1765
rect -31 -1777 2 -1773
rect -39 -1785 2 -1781
rect -47 -1793 2 -1789
rect -55 -1801 2 -1797
rect -62 -1809 2 -1805
rect -69 -1817 2 -1813
rect 2256 -2006 2550 -2002
rect 2256 -2016 2550 -2012
rect 2256 -2025 2550 -2021
rect 2256 -2034 2550 -2030
rect -110 -2039 33 -2035
rect 2256 -2042 2550 -2038
rect 2256 -2050 2550 -2046
rect 2256 -2058 2550 -2054
rect 2256 -2066 2550 -2062
rect 2264 -2105 2309 -2101
rect 2266 -2170 2505 -2166
rect 2266 -2179 2497 -2175
rect 2266 -2188 2489 -2184
rect 2266 -2196 2481 -2192
rect 2266 -2204 2473 -2200
rect 2266 -2212 2465 -2208
rect 2266 -2220 2457 -2216
rect 2266 -2228 2449 -2224
rect -274 -2295 32 -2291
rect -201 -2426 33 -2422
rect 2263 -2493 2404 -2489
rect 2263 -2501 2396 -2497
rect 2263 -2509 2388 -2505
rect 2263 -2517 2380 -2513
rect 2263 -2525 2372 -2521
rect 2263 -2533 2364 -2529
rect 2263 -2542 2356 -2538
rect 2263 -2551 2348 -2547
rect -15 -2919 6 -2915
rect -23 -2928 6 -2924
rect -31 -2936 6 -2932
rect -39 -2944 6 -2940
rect -47 -2952 6 -2948
rect -55 -2960 6 -2956
rect -62 -2968 6 -2964
rect -69 -2976 6 -2972
rect 2262 -3165 2550 -3161
rect 2262 -3175 2550 -3171
rect 2262 -3184 2550 -3180
rect 2262 -3193 2550 -3189
rect -118 -3198 33 -3194
rect 2262 -3201 2550 -3197
rect 2262 -3209 2550 -3205
rect 2262 -3217 2550 -3213
rect 2262 -3225 2550 -3221
rect 2264 -3264 2309 -3260
rect 2266 -3329 2505 -3325
rect 2266 -3338 2497 -3334
rect 2266 -3347 2489 -3343
rect 2266 -3355 2481 -3351
rect 2266 -3363 2473 -3359
rect 2266 -3371 2465 -3367
rect 2266 -3379 2457 -3375
rect 2266 -3387 2449 -3383
rect -282 -3454 33 -3450
rect -209 -3582 33 -3578
rect 2263 -3649 2404 -3645
rect 2263 -3657 2396 -3653
rect 2263 -3665 2388 -3661
rect 2263 -3673 2380 -3669
rect 2263 -3681 2372 -3677
rect 2263 -3689 2364 -3685
rect 2263 -3698 2356 -3694
rect 2263 -3707 2348 -3703
rect -15 -4075 0 -4071
rect -23 -4084 0 -4080
rect -31 -4092 0 -4088
rect -39 -4100 0 -4096
rect -47 -4108 0 -4104
rect -55 -4116 0 -4112
rect -62 -4124 0 -4120
rect -69 -4132 0 -4128
rect 2259 -4321 2550 -4317
rect 2259 -4331 2550 -4327
rect 2259 -4340 2550 -4336
rect 2259 -4349 2550 -4345
rect -126 -4354 33 -4350
rect 2259 -4357 2550 -4353
rect 2259 -4365 2550 -4361
rect 2259 -4373 2550 -4369
rect 2259 -4381 2550 -4377
rect 2264 -4420 2309 -4416
rect 2266 -4485 2505 -4481
rect 2266 -4494 2497 -4490
rect 2266 -4503 2489 -4499
rect 2266 -4511 2481 -4507
rect 2266 -4519 2473 -4515
rect 2266 -4527 2465 -4523
rect 2266 -4535 2457 -4531
rect 2266 -4543 2449 -4539
rect -290 -4610 29 -4606
rect -216 -4740 30 -4736
rect 2263 -4807 2404 -4803
rect 2263 -4815 2396 -4811
rect 2263 -4823 2388 -4819
rect 2263 -4831 2380 -4827
rect 2263 -4839 2372 -4835
rect 2263 -4847 2364 -4843
rect 2263 -4856 2356 -4852
rect 2263 -4865 2348 -4861
rect -15 -5233 0 -5229
rect -23 -5242 0 -5238
rect -31 -5250 0 -5246
rect -39 -5258 0 -5254
rect -47 -5266 0 -5262
rect -55 -5274 0 -5270
rect -62 -5282 1 -5278
rect -69 -5290 14 -5286
rect 2258 -5479 2550 -5475
rect 2258 -5489 2550 -5485
rect 2258 -5498 2550 -5494
rect 2258 -5507 2550 -5503
rect -134 -5512 27 -5508
rect 2258 -5515 2550 -5511
rect 2258 -5523 2550 -5519
rect 2258 -5531 2550 -5527
rect 2258 -5539 2550 -5535
rect 2264 -5578 2309 -5574
rect 2266 -5643 2505 -5639
rect 2266 -5652 2497 -5648
rect 2266 -5661 2489 -5657
rect 2266 -5669 2481 -5665
rect 2266 -5677 2473 -5673
rect 2266 -5685 2465 -5681
rect 2266 -5693 2457 -5689
rect 2266 -5701 2449 -5697
rect -297 -5768 29 -5764
rect -223 -5907 30 -5903
rect 2263 -5974 2404 -5970
rect 2263 -5982 2396 -5978
rect 2263 -5990 2388 -5986
rect 2263 -5998 2380 -5994
rect 2263 -6006 2372 -6002
rect 2263 -6014 2364 -6010
rect 2263 -6023 2356 -6019
rect 2263 -6032 2348 -6028
rect 2260 -6223 2550 -6219
rect 2260 -6233 2550 -6229
rect 2260 -6242 2550 -6238
rect 2260 -6251 2550 -6247
rect 2260 -6259 2550 -6255
rect 2260 -6267 2550 -6263
rect 2260 -6275 2550 -6271
rect 2260 -6283 2550 -6279
rect 2266 -6387 2505 -6383
rect 2266 -6396 2497 -6392
rect 2266 -6405 2489 -6401
rect 2266 -6413 2481 -6409
rect 2266 -6421 2473 -6417
rect 2266 -6429 2465 -6425
rect 2266 -6437 2457 -6433
rect 2266 -6445 2449 -6441
rect -304 -6512 29 -6508
<< m2contact >>
rect 697 2408 701 2412
rect 638 2324 642 2328
rect -521 2301 -517 2305
rect -19 2301 -15 2305
rect -457 2293 -453 2297
rect -27 2293 -23 2297
rect -393 2285 -389 2289
rect -35 2285 -31 2289
rect -329 2277 -325 2281
rect -43 2277 -39 2281
rect -265 2269 -261 2273
rect -51 2269 -47 2273
rect -201 2261 -197 2265
rect -59 2261 -55 2265
rect -137 2253 -133 2257
rect -66 2253 -62 2257
rect -554 2236 -550 2240
rect -490 2228 -486 2232
rect -9 2225 -5 2229
rect -426 2220 -422 2224
rect -362 2212 -358 2216
rect -298 2204 -294 2208
rect -234 2196 -230 2200
rect -170 2188 -166 2192
rect -106 2179 -102 2183
rect -529 2155 -525 2159
rect 2404 2158 2408 2162
rect -465 2147 -461 2151
rect 2396 2150 2400 2154
rect -401 2139 -397 2143
rect 2388 2142 2392 2146
rect -337 2131 -333 2135
rect 2380 2134 2384 2138
rect -273 2123 -269 2127
rect 2372 2126 2376 2130
rect -209 2115 -205 2119
rect 2364 2118 2368 2122
rect -145 2107 -141 2111
rect 2356 2109 2360 2113
rect -81 2099 -77 2103
rect 2348 2100 2352 2104
rect -173 1911 -169 1915
rect -9 1911 -5 1915
rect -19 1732 -15 1736
rect -27 1723 -23 1727
rect -35 1715 -31 1719
rect -43 1707 -39 1711
rect -51 1699 -47 1703
rect -59 1691 -55 1695
rect -66 1683 -62 1687
rect -73 1675 -69 1679
rect -204 1670 -200 1674
rect -204 1617 -200 1621
rect 112 1617 116 1621
rect 13 1586 17 1590
rect -751 1514 -747 1518
rect -735 1506 -731 1510
rect -719 1498 -715 1502
rect -767 1490 -763 1494
rect -367 1453 -363 1457
rect -351 1445 -347 1449
rect -99 1445 -95 1449
rect -335 1437 -331 1441
rect -106 1437 -102 1441
rect -319 1429 -315 1433
rect -114 1429 -110 1433
rect -303 1421 -299 1425
rect -122 1421 -118 1425
rect -287 1413 -283 1417
rect -130 1413 -126 1417
rect -271 1405 -267 1409
rect -138 1405 -134 1409
rect 2309 1387 2313 1391
rect -271 1325 -267 1329
rect 697 1325 701 1329
rect 2505 1322 2509 1326
rect 2497 1313 2501 1317
rect 2489 1304 2493 1308
rect 2481 1296 2485 1300
rect 2473 1288 2477 1292
rect 2465 1280 2469 1284
rect 2457 1272 2461 1276
rect 2449 1264 2453 1268
rect -271 1252 -267 1256
rect 13 1241 17 1245
rect -254 1197 -250 1201
rect -676 1168 -672 1172
rect 13 1168 17 1172
rect -676 1156 -672 1160
rect -666 1156 -662 1160
rect -650 1096 -646 1100
rect -634 1088 -630 1092
rect -569 1087 -565 1091
rect -173 1087 -169 1091
rect -618 1080 -614 1084
rect -528 1079 -524 1083
rect -487 1071 -483 1075
rect -189 1071 -185 1075
rect -446 1063 -442 1067
rect -197 1063 -193 1067
rect -405 1055 -401 1059
rect -205 1055 -201 1059
rect -364 1047 -360 1051
rect -213 1047 -209 1051
rect -323 1039 -319 1043
rect -220 1039 -216 1043
rect -282 1031 -278 1035
rect -227 1031 -223 1035
rect 2404 1012 2408 1016
rect 2396 1004 2400 1008
rect 2388 996 2392 1000
rect 2380 988 2384 992
rect 2372 980 2376 984
rect 2364 972 2368 976
rect 2356 963 2360 967
rect 2348 954 2352 958
rect -19 586 -15 590
rect -27 577 -23 581
rect -35 569 -31 573
rect -43 561 -39 565
rect -51 553 -47 557
rect -59 545 -55 549
rect -66 537 -62 541
rect -73 529 -69 533
rect -99 307 -95 311
rect 112 242 116 246
rect 2309 241 2313 245
rect 2505 176 2509 180
rect 2497 167 2501 171
rect -702 158 -698 162
rect 638 158 642 162
rect 2489 158 2493 162
rect 2481 150 2485 154
rect -702 146 -698 150
rect -692 146 -688 150
rect 2473 142 2477 146
rect 2465 134 2469 138
rect 2457 126 2461 130
rect 2449 118 2453 122
rect -676 70 -672 74
rect -660 62 -656 66
rect -595 59 -591 63
rect -254 59 -250 63
rect -644 54 -640 58
rect -554 51 -550 55
rect -513 43 -509 47
rect -270 43 -266 47
rect -472 35 -468 39
rect -278 35 -274 39
rect -431 27 -427 31
rect -286 27 -282 31
rect -390 19 -386 23
rect -294 19 -290 23
rect -349 11 -345 15
rect -301 11 -297 15
rect -189 -95 -185 -91
rect 2404 -162 2408 -158
rect 2396 -170 2400 -166
rect 2388 -178 2392 -174
rect 2380 -186 2384 -182
rect 2372 -194 2376 -190
rect 2364 -202 2368 -198
rect 2356 -211 2360 -207
rect 2348 -220 2352 -216
rect -19 -588 -15 -584
rect -27 -597 -23 -593
rect -35 -605 -31 -601
rect -43 -613 -39 -609
rect -51 -621 -47 -617
rect -59 -629 -55 -625
rect -66 -637 -62 -633
rect -73 -645 -69 -641
rect -106 -867 -102 -863
rect 2309 -933 2313 -929
rect 2505 -998 2509 -994
rect 2497 -1007 2501 -1003
rect 2489 -1016 2493 -1012
rect 2481 -1024 2485 -1020
rect 2473 -1032 2477 -1028
rect 2465 -1040 2469 -1036
rect 2457 -1048 2461 -1044
rect 2449 -1056 2453 -1052
rect -270 -1123 -266 -1119
rect -197 -1267 -193 -1263
rect 2404 -1334 2408 -1330
rect 2396 -1342 2400 -1338
rect 2388 -1350 2392 -1346
rect 2380 -1358 2384 -1354
rect 2372 -1366 2376 -1362
rect 2364 -1374 2368 -1370
rect 2356 -1383 2360 -1379
rect 2348 -1392 2352 -1388
rect -19 -1760 -15 -1756
rect -27 -1769 -23 -1765
rect -35 -1777 -31 -1773
rect -43 -1785 -39 -1781
rect -51 -1793 -47 -1789
rect -59 -1801 -55 -1797
rect -66 -1809 -62 -1805
rect -73 -1817 -69 -1813
rect -114 -2039 -110 -2035
rect 2309 -2105 2313 -2101
rect 2505 -2170 2509 -2166
rect 2497 -2179 2501 -2175
rect 2489 -2188 2493 -2184
rect 2481 -2196 2485 -2192
rect 2473 -2204 2477 -2200
rect 2465 -2212 2469 -2208
rect 2457 -2220 2461 -2216
rect 2449 -2228 2453 -2224
rect -278 -2295 -274 -2291
rect -205 -2426 -201 -2422
rect 2404 -2493 2408 -2489
rect 2396 -2501 2400 -2497
rect 2388 -2509 2392 -2505
rect 2380 -2517 2384 -2513
rect 2372 -2525 2376 -2521
rect 2364 -2533 2368 -2529
rect 2356 -2542 2360 -2538
rect 2348 -2551 2352 -2547
rect -19 -2919 -15 -2915
rect -27 -2928 -23 -2924
rect -35 -2936 -31 -2932
rect -43 -2944 -39 -2940
rect -51 -2952 -47 -2948
rect -59 -2960 -55 -2956
rect -66 -2968 -62 -2964
rect -73 -2976 -69 -2972
rect -122 -3198 -118 -3194
rect 2309 -3264 2313 -3260
rect 2505 -3329 2509 -3325
rect 2497 -3338 2501 -3334
rect 2489 -3347 2493 -3343
rect 2481 -3355 2485 -3351
rect 2473 -3363 2477 -3359
rect 2465 -3371 2469 -3367
rect 2457 -3379 2461 -3375
rect 2449 -3387 2453 -3383
rect -286 -3454 -282 -3450
rect -213 -3582 -209 -3578
rect 2404 -3649 2408 -3645
rect 2396 -3657 2400 -3653
rect 2388 -3665 2392 -3661
rect 2380 -3673 2384 -3669
rect 2372 -3681 2376 -3677
rect 2364 -3689 2368 -3685
rect 2356 -3698 2360 -3694
rect 2348 -3707 2352 -3703
rect -19 -4075 -15 -4071
rect -27 -4084 -23 -4080
rect -35 -4092 -31 -4088
rect -43 -4100 -39 -4096
rect -51 -4108 -47 -4104
rect -59 -4116 -55 -4112
rect -66 -4124 -62 -4120
rect -73 -4132 -69 -4128
rect -130 -4354 -126 -4350
rect 2309 -4420 2313 -4416
rect 2505 -4485 2509 -4481
rect 2497 -4494 2501 -4490
rect 2489 -4503 2493 -4499
rect 2481 -4511 2485 -4507
rect 2473 -4519 2477 -4515
rect 2465 -4527 2469 -4523
rect 2457 -4535 2461 -4531
rect 2449 -4543 2453 -4539
rect -294 -4610 -290 -4606
rect -220 -4740 -216 -4736
rect 2404 -4807 2408 -4803
rect 2396 -4815 2400 -4811
rect 2388 -4823 2392 -4819
rect 2380 -4831 2384 -4827
rect 2372 -4839 2376 -4835
rect 2364 -4847 2368 -4843
rect 2356 -4856 2360 -4852
rect 2348 -4865 2352 -4861
rect -19 -5233 -15 -5229
rect -27 -5242 -23 -5238
rect -35 -5250 -31 -5246
rect -43 -5258 -39 -5254
rect -51 -5266 -47 -5262
rect -59 -5274 -55 -5270
rect -66 -5282 -62 -5278
rect -73 -5290 -69 -5286
rect -138 -5512 -134 -5508
rect 2309 -5578 2313 -5574
rect 2505 -5643 2509 -5639
rect 2497 -5652 2501 -5648
rect 2489 -5661 2493 -5657
rect 2481 -5669 2485 -5665
rect 2473 -5677 2477 -5673
rect 2465 -5685 2469 -5681
rect 2457 -5693 2461 -5689
rect 2449 -5701 2453 -5697
rect -301 -5768 -297 -5764
rect -227 -5907 -223 -5903
rect 2404 -5974 2408 -5970
rect 2396 -5982 2400 -5978
rect 2388 -5990 2392 -5986
rect 2380 -5998 2384 -5994
rect 2372 -6006 2376 -6002
rect 2364 -6014 2368 -6010
rect 2356 -6023 2360 -6019
rect 2348 -6032 2352 -6028
rect 2505 -6387 2509 -6383
rect 2497 -6396 2501 -6392
rect 2489 -6405 2493 -6401
rect 2481 -6413 2485 -6409
rect 2473 -6421 2477 -6417
rect 2465 -6429 2469 -6425
rect 2457 -6437 2461 -6433
rect 2449 -6445 2453 -6441
rect -308 -6512 -304 -6508
<< metal2 >>
rect -554 2240 -550 2364
rect -529 2159 -525 2364
rect -521 2305 -517 2308
rect -490 2232 -486 2364
rect -465 2151 -461 2364
rect -457 2297 -453 2308
rect -426 2224 -422 2364
rect -401 2143 -397 2364
rect -393 2289 -389 2308
rect -362 2216 -358 2364
rect -337 2135 -333 2364
rect -329 2281 -325 2308
rect -298 2208 -294 2364
rect -273 2127 -269 2364
rect -265 2273 -261 2308
rect -234 2200 -230 2364
rect -209 2119 -205 2364
rect -201 2265 -197 2308
rect -170 2192 -166 2364
rect -145 2111 -141 2364
rect -137 2257 -133 2308
rect -106 2183 -102 2364
rect -81 2103 -77 2364
rect -204 1621 -200 1670
rect -767 1494 -763 1579
rect -751 1518 -747 1571
rect -735 1510 -731 1555
rect -719 1502 -715 1540
rect -367 1457 -363 1579
rect -351 1449 -347 1579
rect -335 1441 -331 1579
rect -319 1433 -315 1579
rect -303 1425 -299 1579
rect -287 1417 -283 1579
rect -271 1409 -267 1579
rect -271 1256 -267 1325
rect -676 1160 -672 1168
rect -650 1100 -646 1152
rect -634 1092 -630 1136
rect -618 1084 -614 1120
rect -569 1091 -565 1105
rect -528 1083 -524 1105
rect -487 1075 -483 1105
rect -446 1067 -442 1105
rect -405 1059 -401 1105
rect -364 1051 -360 1106
rect -323 1043 -319 1105
rect -282 1035 -278 1105
rect -702 150 -698 158
rect -676 74 -672 142
rect -660 66 -656 126
rect -644 58 -640 110
rect -595 63 -591 96
rect -554 55 -550 96
rect -513 47 -509 96
rect -472 39 -468 96
rect -431 31 -427 96
rect -390 23 -386 97
rect -349 15 -345 95
rect -308 -6508 -304 96
rect -254 63 -250 1197
rect -173 1091 -169 1911
rect -73 1679 -69 2308
rect -301 -5764 -297 11
rect -294 -4606 -290 19
rect -286 -3450 -282 27
rect -278 -2291 -274 35
rect -270 -1119 -266 43
rect -227 -5903 -223 1031
rect -220 -4736 -216 1039
rect -213 -3578 -209 1047
rect -205 -2422 -201 1055
rect -197 -1263 -193 1063
rect -189 -91 -185 1071
rect -138 -5508 -134 1405
rect -130 -4350 -126 1413
rect -122 -3194 -118 1421
rect -114 -2035 -110 1429
rect -106 -863 -102 1437
rect -99 311 -95 1445
rect -73 533 -69 1675
rect -73 -641 -69 529
rect -73 -1813 -69 -645
rect -73 -2972 -69 -1817
rect -73 -4128 -69 -2976
rect -73 -5286 -69 -4132
rect -66 1687 -62 2253
rect -66 541 -62 1683
rect -66 -633 -62 537
rect -66 -1805 -62 -637
rect -66 -2964 -62 -1809
rect -66 -4120 -62 -2968
rect -66 -5278 -62 -4124
rect -59 1695 -55 2261
rect -59 549 -55 1691
rect -59 -625 -55 545
rect -59 -1797 -55 -629
rect -59 -2956 -55 -1801
rect -59 -4112 -55 -2960
rect -59 -5270 -55 -4116
rect -51 1703 -47 2269
rect -51 557 -47 1699
rect -51 -617 -47 553
rect -51 -1789 -47 -621
rect -51 -2948 -47 -1793
rect -51 -4104 -47 -2952
rect -51 -5262 -47 -4108
rect -43 1711 -39 2277
rect -43 565 -39 1707
rect -43 -609 -39 561
rect -43 -1781 -39 -613
rect -43 -2940 -39 -1785
rect -43 -4096 -39 -2944
rect -43 -5254 -39 -4100
rect -35 1719 -31 2285
rect -35 573 -31 1715
rect -35 -601 -31 569
rect -35 -1773 -31 -605
rect -35 -2932 -31 -1777
rect -35 -4088 -31 -2936
rect -35 -5246 -31 -4092
rect -27 1727 -23 2293
rect -27 581 -23 1723
rect -27 -593 -23 577
rect -27 -1765 -23 -597
rect -27 -2924 -23 -1769
rect -27 -4080 -23 -2928
rect -27 -5238 -23 -4084
rect -19 1736 -15 2301
rect -9 1915 -5 2225
rect 638 2185 642 2324
rect 697 2269 701 2408
rect -19 590 -15 1732
rect 13 1245 17 1586
rect 13 1172 17 1241
rect 638 1039 642 1253
rect 697 1123 701 1157
rect -19 -584 -15 586
rect 112 246 116 334
rect 638 162 642 293
rect 638 -135 642 158
rect 2309 245 2313 1387
rect 697 -51 701 11
rect -19 -1756 -15 -588
rect 2309 -929 2313 241
rect 638 -1307 642 -932
rect 697 -1223 701 -1163
rect -19 -2915 -15 -1760
rect 638 -2466 642 -2050
rect 2309 -2101 2313 -933
rect 697 -2382 701 -2335
rect -19 -4071 -15 -2919
rect 2309 -3260 2313 -2105
rect 638 -3622 642 -3408
rect 697 -3538 701 -3494
rect -19 -5229 -15 -4075
rect 2309 -4416 2313 -3264
rect 638 -4780 642 -4566
rect 697 -4696 701 -4650
rect 2309 -5574 2313 -4420
rect 638 -5947 642 -5724
rect 697 -5864 701 -5808
rect 2309 -6666 2313 -5578
rect 2348 958 2352 2100
rect 2348 -216 2352 954
rect 2348 -1388 2352 -220
rect 2348 -2547 2352 -1392
rect 2348 -3703 2352 -2551
rect 2348 -4861 2352 -3707
rect 2348 -6028 2352 -4865
rect 2348 -6666 2352 -6032
rect 2356 967 2360 2109
rect 2356 -207 2360 963
rect 2356 -1379 2360 -211
rect 2356 -2538 2360 -1383
rect 2356 -3694 2360 -2542
rect 2356 -4852 2360 -3698
rect 2356 -6019 2360 -4856
rect 2356 -6666 2360 -6023
rect 2364 976 2368 2118
rect 2364 -198 2368 972
rect 2364 -1370 2368 -202
rect 2364 -2529 2368 -1374
rect 2364 -3685 2368 -2533
rect 2364 -4843 2368 -3689
rect 2364 -6010 2368 -4847
rect 2364 -6666 2368 -6014
rect 2372 984 2376 2126
rect 2372 -190 2376 980
rect 2372 -1362 2376 -194
rect 2372 -2521 2376 -1366
rect 2372 -3677 2376 -2525
rect 2372 -4835 2376 -3681
rect 2372 -6002 2376 -4839
rect 2372 -6666 2376 -6006
rect 2380 992 2384 2134
rect 2380 -182 2384 988
rect 2380 -1354 2384 -186
rect 2380 -2513 2384 -1358
rect 2380 -3669 2384 -2517
rect 2380 -4827 2384 -3673
rect 2380 -5994 2384 -4831
rect 2380 -6666 2384 -5998
rect 2388 1000 2392 2142
rect 2388 -174 2392 996
rect 2388 -1346 2392 -178
rect 2388 -2505 2392 -1350
rect 2388 -3661 2392 -2509
rect 2388 -4819 2392 -3665
rect 2388 -5986 2392 -4823
rect 2388 -6666 2392 -5990
rect 2396 1008 2400 2150
rect 2396 -166 2400 1004
rect 2396 -1338 2400 -170
rect 2396 -2497 2400 -1342
rect 2396 -3653 2400 -2501
rect 2396 -4811 2400 -3657
rect 2396 -5978 2400 -4815
rect 2396 -6666 2400 -5982
rect 2404 1016 2408 2158
rect 2404 -158 2408 1012
rect 2404 -1330 2408 -162
rect 2404 -2489 2408 -1334
rect 2404 -3645 2408 -2493
rect 2404 -4803 2408 -3649
rect 2404 -5970 2408 -4807
rect 2404 -6666 2408 -5974
rect 2449 122 2453 1264
rect 2449 -1052 2453 118
rect 2449 -2224 2453 -1056
rect 2449 -3383 2453 -2228
rect 2449 -4539 2453 -3387
rect 2449 -5697 2453 -4543
rect 2449 -6441 2453 -5701
rect 2449 -6666 2453 -6445
rect 2457 130 2461 1272
rect 2457 -1044 2461 126
rect 2457 -2216 2461 -1048
rect 2457 -3375 2461 -2220
rect 2457 -4531 2461 -3379
rect 2457 -5689 2461 -4535
rect 2457 -6433 2461 -5693
rect 2457 -6666 2461 -6437
rect 2465 138 2469 1280
rect 2465 -1036 2469 134
rect 2465 -2208 2469 -1040
rect 2465 -3367 2469 -2212
rect 2465 -4523 2469 -3371
rect 2465 -5681 2469 -4527
rect 2465 -6425 2469 -5685
rect 2465 -6666 2469 -6429
rect 2473 146 2477 1288
rect 2473 -1028 2477 142
rect 2473 -2200 2477 -1032
rect 2473 -3359 2477 -2204
rect 2473 -4515 2477 -3363
rect 2473 -5673 2477 -4519
rect 2473 -6417 2477 -5677
rect 2473 -6666 2477 -6421
rect 2481 154 2485 1296
rect 2481 -1020 2485 150
rect 2481 -2192 2485 -1024
rect 2481 -3351 2485 -2196
rect 2481 -4507 2485 -3355
rect 2481 -5665 2485 -4511
rect 2481 -6409 2485 -5669
rect 2481 -6666 2485 -6413
rect 2489 162 2493 1304
rect 2489 -1012 2493 158
rect 2489 -2184 2493 -1016
rect 2489 -3343 2493 -2188
rect 2489 -4499 2493 -3347
rect 2489 -5657 2493 -4503
rect 2489 -6401 2493 -5661
rect 2489 -6666 2493 -6405
rect 2497 171 2501 1313
rect 2497 -1003 2501 167
rect 2497 -2175 2501 -1007
rect 2497 -3334 2501 -2179
rect 2497 -4490 2501 -3338
rect 2497 -5648 2501 -4494
rect 2497 -6392 2501 -5652
rect 2497 -6666 2501 -6396
rect 2505 180 2509 1322
rect 2505 -994 2509 176
rect 2505 -2166 2509 -998
rect 2505 -3325 2509 -2170
rect 2505 -4481 2509 -3329
rect 2505 -5639 2509 -4485
rect 2505 -6383 2509 -5643
rect 2505 -6666 2509 -6387
use REG0  REG0_0
timestamp 1746042099
transform 1 0 -1 0 1 -6554
box 30 -2 2267 696
use REG8  REG8_6
timestamp 1746070328
transform 1 0 29 0 1 -5443
box -29 -376 2237 759
use REG8  REG8_5
timestamp 1746070328
transform 1 0 29 0 1 -4285
box -29 -376 2237 759
use REG8  REG8_4
timestamp 1746070328
transform 1 0 29 0 1 -3129
box -29 -376 2237 759
use REG8  REG8_3
timestamp 1746070328
transform 1 0 29 0 1 -1970
box -29 -376 2237 759
use REG8  REG8_2
timestamp 1746070328
transform 1 0 29 0 1 -798
box -29 -376 2237 759
use Decoder_4x8  Decoder_4x8_1
timestamp 1742681920
transform 1 0 -634 0 1 158
box -64 -64 336 95
use REG8  REG8_1
timestamp 1746070328
transform 1 0 29 0 1 376
box -29 -376 2237 759
use Decoder_4x8  Decoder_4x8_0
timestamp 1742681920
transform 1 0 -608 0 1 1168
box -64 -64 336 95
use REG8  REG8_7
timestamp 1746070328
transform 1 0 29 0 1 1522
box -29 -376 2237 759
use 8bitMUX2to1  8bitMUX2to1_0
timestamp 1746042099
transform 1 0 -583 0 1 2308
box 0 0 520 107
use Decoder_Inv_4x8  Decoder_Inv_4x8_0
timestamp 1743018986
transform 1 0 -773 0 1 1522
box 0 -56 528 159
<< labels >>
rlabel metal2 2311 -6664 2311 -6664 1 CLK
rlabel metal2 2406 -6664 2406 -6664 1 B0
rlabel metal2 2398 -6664 2398 -6664 1 B1
rlabel metal2 2390 -6664 2390 -6664 1 B2
rlabel metal2 2382 -6664 2382 -6664 1 B3
rlabel metal2 2374 -6664 2374 -6664 1 B4
rlabel metal2 2366 -6664 2366 -6664 1 B5
rlabel metal2 2358 -6664 2358 -6664 1 B6
rlabel metal2 2350 -6664 2350 -6664 1 B7
rlabel metal2 2507 -6664 2507 -6664 1 A0
rlabel metal2 2499 -6664 2499 -6664 1 A1
rlabel metal2 2491 -6664 2491 -6664 1 A2
rlabel metal2 2483 -6664 2483 -6664 1 A3
rlabel metal2 2475 -6664 2475 -6664 1 A4
rlabel metal2 2467 -6664 2467 -6664 1 A5
rlabel metal2 2459 -6664 2459 -6664 1 A6
rlabel metal2 2451 -6664 2451 -6664 1 A7
rlabel metal1 -808 2238 -808 2238 1 C0
rlabel metal1 -808 2230 -808 2230 1 C1
rlabel metal1 -808 2222 -808 2222 1 C2
rlabel metal1 -808 2214 -808 2214 1 C3
rlabel metal1 -808 2206 -808 2206 1 C4
rlabel metal1 -808 2198 -808 2198 1 C5
rlabel metal1 -808 2190 -808 2190 1 C6
rlabel metal1 -808 2181 -808 2181 1 C7
rlabel metal1 -808 2157 -808 2157 1 Imm0
rlabel metal1 -808 2149 -808 2149 1 Imm1
rlabel metal1 -808 2141 -808 2141 1 Imm2
rlabel metal1 -808 2133 -808 2133 1 Imm3
rlabel metal1 -808 2125 -808 2125 1 Imm4
rlabel metal1 -808 2117 -808 2117 1 Imm5
rlabel metal1 -808 2109 -808 2109 1 Imm6
rlabel metal1 -808 2101 -808 2101 1 Imm7
rlabel metal1 217 2410 217 2410 1 VDD
rlabel metal1 218 2326 218 2326 1 VSS
rlabel metal1 -808 72 -808 72 1 A_sel0
rlabel metal1 -808 64 -808 64 1 A_sel1
rlabel metal1 -808 56 -808 56 1 A_sel2
rlabel metal1 -808 1098 -808 1098 1 B_sel0
rlabel metal1 -808 1090 -808 1090 1 B_sel1
rlabel metal1 -808 1082 -808 1082 1 B_sel2
rlabel metal1 -808 1516 -808 1516 1 C_sel0
rlabel metal1 -808 1508 -808 1508 1 C_sel1
rlabel metal1 -808 1500 -808 1500 1 C_sel2
rlabel metal1 -808 1492 -808 1492 1 C_sel3
rlabel metal1 -808 2370 -808 2370 1 Imm_en
rlabel metal1 2548 1488 2548 1488 1 reg_zero0
rlabel metal1 2548 1478 2548 1478 1 reg_zero1
rlabel metal1 2548 1469 2548 1469 1 reg_zero2
rlabel metal1 2547 1460 2547 1460 1 reg_zero3
rlabel metal1 2545 1452 2545 1452 1 reg_zero4
rlabel metal1 2545 1444 2545 1444 1 reg_zero5
rlabel metal1 2545 1436 2545 1436 1 reg_zero6
rlabel metal1 2546 1428 2546 1428 1 reg_zero7
rlabel metal2 -17 1741 -17 1741 1 check
rlabel metal1 2548 342 2548 342 1 reg_one0
rlabel metal1 2548 332 2548 332 1 reg_one1
rlabel metal1 2548 323 2548 323 1 reg_one2
rlabel metal1 2548 314 2548 314 1 reg_one3
rlabel metal1 2548 306 2548 306 1 reg_one4
rlabel metal1 2548 298 2548 298 1 reg_one5
rlabel metal1 2548 290 2548 290 1 reg_one6
rlabel metal1 2548 282 2548 282 1 reg_one7
rlabel metal1 2547 -832 2547 -832 1 reg_two0
rlabel metal1 2547 -842 2547 -842 1 reg_two1
rlabel metal1 2547 -851 2547 -851 1 reg_two2
rlabel metal1 2547 -860 2547 -860 1 reg_two3
rlabel metal1 2547 -868 2547 -868 1 reg_two4
rlabel metal1 2547 -876 2547 -876 1 reg_two5
rlabel metal1 2547 -884 2547 -884 1 reg_two6
rlabel metal1 2547 -892 2547 -892 1 reg_two7
rlabel metal1 2546 -2004 2546 -2004 1 reg_three0
rlabel metal1 2546 -2014 2546 -2014 1 reg_three1
rlabel metal1 2547 -2023 2547 -2023 1 reg_three2
rlabel metal1 2547 -2032 2547 -2032 1 reg_three3
rlabel metal1 2547 -2040 2547 -2040 1 reg_three4
rlabel metal1 2547 -2048 2547 -2048 1 reg_three5
rlabel metal1 2547 -2056 2547 -2056 1 reg_three6
rlabel metal1 2547 -2064 2547 -2064 1 reg_three7
rlabel metal1 2546 -3163 2546 -3163 1 reg_four0
rlabel metal1 2547 -3173 2547 -3173 1 reg_four1
rlabel metal1 2547 -3182 2547 -3182 1 reg_four2
rlabel metal1 2547 -3191 2547 -3191 1 reg_four3
rlabel metal1 2547 -3199 2547 -3199 1 reg_four4
rlabel metal1 2547 -3207 2547 -3207 1 reg_four5
rlabel metal1 2547 -3215 2547 -3215 1 reg_four6
rlabel metal1 2547 -3223 2547 -3223 1 reg_four7
rlabel metal1 2547 -4319 2547 -4319 1 reg_five0
rlabel metal1 2547 -4329 2547 -4329 1 reg_five1
rlabel metal1 2547 -4338 2547 -4338 1 reg_five2
rlabel metal1 2547 -4347 2547 -4347 1 reg_five3
rlabel metal1 2547 -4355 2547 -4355 1 reg_five4
rlabel metal1 2547 -4363 2547 -4363 1 reg_five5
rlabel metal1 2547 -4371 2547 -4371 1 reg_five6
rlabel metal1 2547 -4379 2547 -4379 1 reg_five7
rlabel metal1 2547 -5477 2547 -5477 1 reg_six0
rlabel metal1 2547 -5487 2547 -5487 1 reg_six1
rlabel metal1 2547 -5496 2547 -5496 1 reg_six2
rlabel metal1 2547 -5505 2547 -5505 1 reg_six3
rlabel metal1 2546 -5513 2546 -5513 1 reg_six4
rlabel metal1 2546 -5521 2546 -5521 1 reg_six5
rlabel metal1 2546 -5529 2546 -5529 1 reg_six6
rlabel metal1 2547 -5537 2547 -5537 1 reg_six7
rlabel metal1 2546 -6221 2546 -6221 1 reg_seven0
rlabel metal1 2546 -6231 2546 -6231 1 reg_seven1
rlabel metal1 2546 -6240 2546 -6240 1 reg_seven2
rlabel metal1 2546 -6249 2546 -6249 1 reg_seven3
rlabel metal1 2546 -6257 2546 -6257 1 reg_seven4
rlabel metal1 2546 -6265 2546 -6265 1 reg_seven5
rlabel metal1 2546 -6273 2546 -6273 1 reg_seven6
rlabel metal1 2546 -6281 2546 -6281 1 reg_seven7
<< end >>
