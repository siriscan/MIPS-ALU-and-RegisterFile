magic
tech scmos
timestamp 1746750801
<< nwell >>
rect -44 1784 -18 1788
rect -407 1521 -372 1529
rect -407 1517 -401 1521
rect -182 600 -178 604
rect -132 600 -128 604
rect 100 600 3465 604
<< polysilicon >>
rect 728 1741 730 1744
<< metal1 >>
rect -46 1784 -18 1788
rect 731 1742 735 1743
rect 704 1737 708 1741
rect -37 1725 -33 1729
rect 731 1716 735 1724
rect -413 1709 -407 1713
rect -403 1709 -50 1713
rect -413 1700 -330 1704
rect -326 1700 -40 1704
rect -411 1692 -294 1696
rect -290 1692 6 1696
rect -411 1684 -382 1688
rect -378 1684 -37 1688
rect 2335 1684 3745 1688
rect -411 1676 -398 1680
rect -394 1676 -29 1680
rect 636 1676 639 1680
rect 2335 1676 3685 1680
rect 3689 1676 3745 1680
rect 637 1669 641 1673
rect 2335 1668 3693 1672
rect 3697 1668 3745 1672
rect 2335 1660 3701 1664
rect 3705 1660 3745 1664
rect -2 1653 6 1657
rect 2335 1652 3709 1656
rect 3713 1652 3745 1656
rect -417 1645 -122 1649
rect -118 1645 6 1649
rect 2335 1644 3717 1648
rect 3721 1644 3745 1648
rect -417 1637 -114 1641
rect -110 1637 6 1641
rect 2335 1636 3725 1640
rect 3729 1636 3745 1640
rect -417 1629 -106 1633
rect -102 1629 6 1633
rect 2335 1628 3733 1632
rect 3737 1628 3745 1632
rect -417 1621 -98 1625
rect -94 1621 6 1625
rect 2335 1620 3741 1624
rect -417 1613 -90 1617
rect -86 1613 6 1617
rect -417 1605 -82 1609
rect -78 1605 6 1609
rect -417 1597 -74 1601
rect -70 1597 6 1601
rect -417 1589 -66 1593
rect -62 1589 6 1593
rect -417 1581 -58 1585
rect -54 1581 6 1585
rect -417 1573 -50 1577
rect -46 1573 6 1577
rect -417 1565 -42 1569
rect -38 1565 6 1569
rect -417 1557 -34 1561
rect -30 1557 6 1561
rect -417 1549 -26 1553
rect -22 1549 6 1553
rect -417 1541 -18 1545
rect -14 1541 6 1545
rect -417 1533 -10 1537
rect -6 1533 6 1537
rect -417 1525 -2 1529
rect 2 1525 6 1529
rect -403 1517 -398 1521
rect -132 1517 5 1521
rect -382 1477 -378 1486
rect -314 1473 -310 1477
rect -382 1452 -378 1463
rect -132 1433 5 1437
rect -126 1425 7 1429
rect -118 1417 7 1421
rect 541 1417 3685 1421
rect 3689 1417 3745 1421
rect -110 1409 7 1413
rect 541 1409 3693 1413
rect 3697 1409 3745 1413
rect -394 1401 -278 1405
rect -102 1401 7 1405
rect 541 1401 3701 1405
rect 3705 1401 3745 1405
rect -94 1393 7 1397
rect 541 1393 3709 1397
rect 3713 1393 3745 1397
rect -233 1385 -130 1389
rect -86 1385 7 1389
rect 541 1385 3717 1389
rect 3721 1385 3745 1389
rect -78 1377 7 1381
rect 541 1377 3725 1381
rect 3729 1377 3745 1381
rect -70 1369 7 1373
rect 541 1369 3733 1373
rect 3737 1369 3745 1373
rect -62 1361 7 1365
rect 541 1361 3741 1365
rect -54 1354 7 1358
rect -46 1346 7 1350
rect -38 1338 7 1342
rect -30 1330 7 1334
rect -22 1322 7 1326
rect -14 1314 7 1318
rect -6 1306 7 1310
rect 2 1298 7 1302
rect -403 1290 4 1294
rect -326 1206 4 1210
rect -200 1198 4 1202
rect -118 1190 5 1194
rect 572 1190 3685 1194
rect 3689 1190 3745 1194
rect -110 1182 5 1186
rect 572 1182 3693 1186
rect 3697 1182 3745 1186
rect -102 1174 6 1178
rect 572 1174 3701 1178
rect 3705 1174 3745 1178
rect -94 1166 6 1170
rect 572 1166 3709 1170
rect 3713 1166 3745 1170
rect -86 1158 6 1162
rect 572 1158 3717 1162
rect 3721 1158 3745 1162
rect -78 1150 6 1154
rect 572 1150 3725 1154
rect 3729 1150 3745 1154
rect -70 1142 6 1146
rect 572 1142 3733 1146
rect 3737 1142 3745 1146
rect -62 1134 6 1138
rect 572 1134 3741 1138
rect -54 1126 6 1130
rect -46 1118 6 1122
rect -38 1110 6 1114
rect -30 1102 6 1106
rect -22 1094 6 1098
rect -14 1086 6 1090
rect -6 1078 4 1082
rect 2 1070 4 1074
rect -403 1060 4 1064
rect -326 976 4 980
rect -167 968 6 972
rect -118 956 6 960
rect 796 956 3685 960
rect 3689 956 3745 960
rect -110 948 6 952
rect 796 948 3693 952
rect 3697 948 3745 952
rect -102 940 6 944
rect 796 940 3701 944
rect 3705 940 3745 944
rect -94 932 6 936
rect 796 932 3709 936
rect 3713 932 3745 936
rect -86 924 6 928
rect 796 924 3717 928
rect 3721 924 3745 928
rect -78 916 6 920
rect 796 916 3725 920
rect 3729 916 3745 920
rect -70 908 6 912
rect 796 908 3733 912
rect 3737 908 3745 912
rect -62 900 6 904
rect 796 900 3741 904
rect -54 892 6 896
rect -46 884 6 888
rect -38 876 6 880
rect -30 868 6 872
rect -22 860 6 864
rect -14 852 6 856
rect -6 844 6 848
rect 2 836 6 840
rect -403 828 5 832
rect -326 744 4 748
rect -134 736 4 740
rect -118 728 4 732
rect 444 728 3685 732
rect 3689 728 3745 732
rect -110 720 4 724
rect 444 720 3693 724
rect 3697 720 3745 724
rect -102 712 4 716
rect 444 712 3701 716
rect 3705 712 3745 716
rect -94 704 4 708
rect 444 704 3709 708
rect 3713 704 3745 708
rect -86 696 4 700
rect 444 696 3717 700
rect 3721 696 3745 700
rect -78 688 4 692
rect 444 688 3725 692
rect 3729 688 3745 692
rect -70 680 4 684
rect 444 680 3733 684
rect 3737 680 3745 684
rect -62 672 4 676
rect 444 672 3741 676
rect -54 664 4 668
rect -46 656 4 660
rect -38 648 4 652
rect -30 640 4 644
rect -22 632 4 636
rect -14 624 4 628
rect -6 616 4 620
rect 2 608 4 612
rect -403 600 -178 604
rect -132 600 5 604
rect 100 600 3465 604
rect -290 556 -179 560
rect -167 540 -162 544
rect -326 516 -180 520
rect -132 516 -130 520
rect -126 516 6 520
rect 100 516 3465 520
rect -394 508 -153 512
rect -378 500 -145 504
rect 3679 500 3685 504
rect 3689 500 3745 504
rect -417 492 7 496
rect 3679 492 3693 496
rect 3697 492 3745 496
rect 3678 484 3701 488
rect 3705 484 3745 488
rect -118 476 7 480
rect 3475 476 3479 480
rect 3679 476 3709 480
rect 3713 476 3745 480
rect -110 468 7 472
rect 3475 468 3479 472
rect 3679 468 3680 472
rect 3681 468 3717 472
rect 3721 468 3745 472
rect -102 460 7 464
rect 3475 460 3479 464
rect 3679 460 3680 464
rect 3681 460 3725 464
rect 3729 460 3745 464
rect -94 452 7 456
rect 3475 452 3479 456
rect 3679 452 3680 456
rect 3681 452 3733 456
rect 3737 452 3745 456
rect -86 444 7 448
rect 3475 444 3479 448
rect 3681 444 3741 448
rect -78 436 7 440
rect 3475 436 3479 440
rect -70 428 7 432
rect 3475 428 3479 432
rect -62 420 7 424
rect 3475 420 3479 424
rect -417 404 8 408
rect -54 396 7 400
rect -46 388 7 392
rect -38 380 7 384
rect -134 316 9 320
rect -403 308 -158 312
rect -128 308 4 312
rect -290 282 -140 286
rect -378 265 -148 269
rect -394 248 -157 252
rect -326 224 -159 228
rect -137 224 -133 228
rect -128 224 4 228
rect 2392 208 3685 212
rect 3689 208 3745 212
rect 2392 200 3693 204
rect 3697 200 3745 204
rect 2392 192 3701 196
rect 3705 192 3745 196
rect 2392 184 3709 188
rect 3713 184 3745 188
rect 2392 176 3717 180
rect 3721 176 3745 180
rect 2392 168 3725 172
rect 3729 168 3745 172
rect 2392 160 3733 164
rect 3737 160 3745 164
rect 2392 152 3741 156
rect -118 136 6 140
rect -110 128 6 132
rect -102 120 6 124
rect -94 112 6 116
rect -86 104 6 108
rect -78 96 6 100
rect -70 88 6 92
rect -62 80 6 84
rect -54 72 6 76
rect -46 64 6 68
rect -38 56 6 60
rect -30 48 6 52
rect -22 40 6 44
rect -14 32 6 36
rect -6 24 6 28
rect 2 16 6 20
rect -129 8 6 12
<< m2contact >>
rect -50 1784 -46 1788
rect -29 1747 -25 1751
rect -37 1729 -33 1733
rect -407 1709 -403 1713
rect -50 1709 -46 1713
rect -6 1712 -2 1716
rect -330 1700 -326 1704
rect -294 1692 -290 1696
rect 6 1692 10 1696
rect -382 1684 -378 1688
rect -37 1684 -33 1688
rect -398 1676 -394 1680
rect -29 1676 -25 1680
rect 3685 1676 3689 1680
rect 3693 1668 3697 1672
rect 3701 1660 3705 1664
rect -6 1653 -2 1657
rect 3709 1652 3713 1656
rect -122 1645 -118 1649
rect 3717 1644 3721 1648
rect -114 1637 -110 1641
rect 3725 1636 3729 1640
rect -106 1629 -102 1633
rect 3733 1628 3737 1632
rect -98 1621 -94 1625
rect 3741 1620 3745 1624
rect -90 1613 -86 1617
rect -82 1605 -78 1609
rect -74 1597 -70 1601
rect -66 1589 -62 1593
rect -58 1581 -54 1585
rect -50 1573 -46 1577
rect -42 1565 -38 1569
rect -34 1557 -30 1561
rect -26 1549 -22 1553
rect -18 1541 -14 1545
rect -10 1533 -6 1537
rect -2 1525 2 1529
rect -407 1517 -403 1521
rect -382 1486 -378 1490
rect -398 1477 -394 1481
rect -382 1448 -378 1452
rect -130 1437 -126 1441
rect -330 1433 -326 1437
rect -130 1425 -126 1429
rect -122 1417 -118 1421
rect 3685 1417 3689 1421
rect -114 1409 -110 1413
rect 3693 1409 3697 1413
rect -398 1401 -394 1405
rect -106 1401 -102 1405
rect 3701 1401 3705 1405
rect -98 1393 -94 1397
rect 3709 1393 3713 1397
rect -237 1385 -233 1389
rect -130 1385 -126 1389
rect -90 1385 -86 1389
rect 3717 1385 3721 1389
rect -82 1377 -78 1381
rect 3725 1377 3729 1381
rect -74 1369 -70 1373
rect 3733 1369 3737 1373
rect -66 1361 -62 1365
rect 3741 1361 3745 1365
rect -58 1354 -54 1358
rect -50 1346 -46 1350
rect -42 1338 -38 1342
rect -34 1330 -30 1334
rect -26 1322 -22 1326
rect -18 1314 -14 1318
rect -10 1306 -6 1310
rect -2 1298 2 1302
rect -407 1290 -403 1294
rect -330 1206 -326 1210
rect -204 1198 -200 1202
rect -122 1190 -118 1194
rect 3685 1190 3689 1194
rect -114 1182 -110 1186
rect 3693 1182 3697 1186
rect -106 1174 -102 1178
rect 3701 1174 3705 1178
rect -98 1166 -94 1170
rect 3709 1166 3713 1170
rect -90 1158 -86 1162
rect 3717 1158 3721 1162
rect -82 1150 -78 1154
rect 3725 1150 3729 1154
rect -74 1142 -70 1146
rect 3733 1142 3737 1146
rect -66 1134 -62 1138
rect 3741 1134 3745 1138
rect -58 1126 -54 1130
rect -50 1118 -46 1122
rect -42 1110 -38 1114
rect -34 1102 -30 1106
rect -26 1094 -22 1098
rect -18 1086 -14 1090
rect -10 1078 -6 1082
rect -2 1070 2 1074
rect -407 1060 -403 1064
rect -330 976 -326 980
rect -171 968 -167 972
rect -122 956 -118 960
rect 3685 956 3689 960
rect -114 948 -110 952
rect 3693 948 3697 952
rect -106 940 -102 944
rect 3701 940 3705 944
rect -98 932 -94 936
rect 3709 932 3713 936
rect -90 924 -86 928
rect 3717 924 3721 928
rect -82 916 -78 920
rect 3725 916 3729 920
rect -74 908 -70 912
rect 3733 908 3737 912
rect -66 900 -62 904
rect 3741 900 3745 904
rect -58 892 -54 896
rect -50 884 -46 888
rect -42 876 -38 880
rect -34 868 -30 872
rect -26 860 -22 864
rect -18 852 -14 856
rect -10 844 -6 848
rect -2 836 2 840
rect -407 828 -403 832
rect -330 744 -326 748
rect -138 736 -134 740
rect -122 728 -118 732
rect 3685 728 3689 732
rect -114 720 -110 724
rect 3693 720 3697 724
rect -106 712 -102 716
rect 3701 712 3705 716
rect -98 704 -94 708
rect 3709 704 3713 708
rect -90 696 -86 700
rect 3717 696 3721 700
rect -82 688 -78 692
rect 3725 688 3729 692
rect -74 680 -70 684
rect 3733 680 3737 684
rect -66 672 -62 676
rect 3741 672 3745 676
rect -58 664 -54 668
rect -50 656 -46 660
rect -42 648 -38 652
rect -34 640 -30 644
rect -26 632 -22 636
rect -18 624 -14 628
rect -10 616 -6 620
rect -2 608 2 612
rect -407 600 -403 604
rect -145 570 -141 574
rect -294 556 -290 560
rect -153 553 -149 557
rect -138 528 -134 532
rect -330 516 -326 520
rect -130 516 -126 520
rect -398 508 -394 512
rect -153 508 -149 512
rect -382 500 -378 504
rect -145 500 -141 504
rect 3685 500 3689 504
rect 3693 492 3697 496
rect 3701 484 3705 488
rect -122 476 -118 480
rect 3709 476 3713 480
rect -114 468 -110 472
rect 3717 468 3721 472
rect -106 460 -102 464
rect 3725 460 3729 464
rect -98 452 -94 456
rect 3733 452 3737 456
rect -90 444 -86 448
rect 3741 444 3745 448
rect -82 436 -78 440
rect -74 428 -70 432
rect -66 420 -62 424
rect -58 396 -54 400
rect -50 388 -46 392
rect -42 380 -38 384
rect -138 316 -134 320
rect -407 308 -403 312
rect -294 282 -290 286
rect -382 265 -378 269
rect -398 248 -394 252
rect -133 236 -129 240
rect -330 224 -326 228
rect 3685 208 3689 212
rect 3693 200 3697 204
rect 3701 192 3705 196
rect 3709 184 3713 188
rect 3717 176 3721 180
rect 3725 168 3729 172
rect 3733 160 3737 164
rect 3741 152 3745 156
rect -122 136 -118 140
rect -114 128 -110 132
rect -106 120 -102 124
rect -98 112 -94 116
rect -90 104 -86 108
rect -82 96 -78 100
rect -74 88 -70 92
rect -66 80 -62 84
rect -58 72 -54 76
rect -50 64 -46 68
rect -42 56 -38 60
rect -34 48 -30 52
rect -26 40 -22 44
rect -18 32 -14 36
rect -10 24 -6 28
rect -2 16 2 20
rect -133 8 -129 12
<< metal2 >>
rect -50 1713 -46 1784
rect -407 1521 -403 1709
rect -407 1294 -403 1517
rect -398 1481 -394 1676
rect -382 1490 -378 1684
rect -407 1064 -403 1290
rect -407 832 -403 1060
rect -407 604 -403 828
rect -407 312 -403 600
rect -398 1405 -394 1456
rect -398 512 -394 1401
rect -398 252 -394 508
rect -382 504 -378 1448
rect -382 269 -378 500
rect -330 1437 -326 1700
rect -294 1473 -290 1692
rect -37 1688 -33 1729
rect -29 1680 -25 1747
rect -6 1657 -2 1712
rect -330 1210 -326 1433
rect -330 980 -326 1206
rect -330 748 -326 976
rect -330 520 -326 744
rect -330 228 -326 516
rect -294 560 -290 1417
rect -130 1389 -126 1425
rect -204 1202 -200 1389
rect -171 972 -167 1389
rect -138 740 -134 1389
rect -122 1421 -118 1645
rect -122 1194 -118 1417
rect -122 960 -118 1190
rect -122 732 -118 956
rect -294 286 -290 556
rect -153 512 -149 553
rect -145 504 -141 570
rect -138 320 -134 528
rect -122 480 -118 728
rect -133 12 -129 236
rect -122 140 -118 476
rect -114 1413 -110 1637
rect -114 1186 -110 1409
rect -114 952 -110 1182
rect -114 724 -110 948
rect -114 472 -110 720
rect -114 132 -110 468
rect -106 1405 -102 1629
rect -106 1178 -102 1401
rect -106 944 -102 1174
rect -106 716 -102 940
rect -106 464 -102 712
rect -106 124 -102 460
rect -98 1397 -94 1621
rect -98 1170 -94 1393
rect -98 936 -94 1166
rect -98 708 -94 932
rect -98 456 -94 704
rect -98 116 -94 452
rect -90 1389 -86 1613
rect -90 1162 -86 1385
rect -90 928 -86 1158
rect -90 700 -86 924
rect -90 448 -86 696
rect -90 108 -86 444
rect -82 1381 -78 1605
rect -82 1154 -78 1377
rect -82 920 -78 1150
rect -82 692 -78 916
rect -82 440 -78 688
rect -82 100 -78 436
rect -74 1373 -70 1597
rect -74 1146 -70 1369
rect -74 912 -70 1142
rect -74 684 -70 908
rect -74 432 -70 680
rect -74 92 -70 428
rect -66 1365 -62 1589
rect -66 1138 -62 1361
rect -66 904 -62 1134
rect -66 676 -62 900
rect -66 424 -62 672
rect -66 84 -62 420
rect -58 1358 -54 1581
rect -58 1130 -54 1354
rect -58 896 -54 1126
rect -58 668 -54 892
rect -58 400 -54 664
rect -58 76 -54 396
rect -50 1350 -46 1573
rect -50 1122 -46 1346
rect -50 888 -46 1118
rect -50 660 -46 884
rect -50 392 -46 656
rect -50 68 -46 388
rect -42 1342 -38 1565
rect -42 1114 -38 1338
rect -42 880 -38 1110
rect -42 652 -38 876
rect -42 384 -38 648
rect -42 60 -38 380
rect -34 1334 -30 1557
rect -34 1106 -30 1330
rect -34 872 -30 1102
rect -34 644 -30 868
rect -34 52 -30 640
rect -26 1326 -22 1549
rect -26 1098 -22 1322
rect -26 864 -22 1094
rect -26 636 -22 860
rect -26 44 -22 632
rect -18 1318 -14 1541
rect -18 1090 -14 1314
rect -18 856 -14 1086
rect -18 628 -14 852
rect -18 36 -14 624
rect -10 1310 -6 1533
rect -10 1082 -6 1306
rect -10 848 -6 1078
rect -10 620 -6 844
rect -10 28 -6 616
rect -2 1302 2 1525
rect -2 1074 2 1298
rect -2 840 2 1070
rect -2 612 2 836
rect -2 20 2 608
rect 3685 1421 3689 1676
rect 3685 1194 3689 1417
rect 3685 960 3689 1190
rect 3685 732 3689 956
rect 3685 504 3689 728
rect 3685 212 3689 500
rect 3693 1413 3697 1668
rect 3693 1186 3697 1409
rect 3693 952 3697 1182
rect 3693 724 3697 948
rect 3693 496 3697 720
rect 3693 204 3697 492
rect 3701 1405 3705 1660
rect 3701 1178 3705 1401
rect 3701 944 3705 1174
rect 3701 716 3705 940
rect 3701 488 3705 712
rect 3701 196 3705 484
rect 3709 1397 3713 1652
rect 3709 1170 3713 1393
rect 3709 936 3713 1166
rect 3709 708 3713 932
rect 3709 480 3713 704
rect 3709 188 3713 476
rect 3717 1389 3721 1644
rect 3717 1162 3721 1385
rect 3717 928 3721 1158
rect 3717 700 3721 924
rect 3717 472 3721 696
rect 3717 180 3721 468
rect 3725 1381 3729 1636
rect 3725 1154 3729 1377
rect 3725 920 3729 1150
rect 3725 692 3729 916
rect 3725 464 3729 688
rect 3725 172 3729 460
rect 3733 1373 3737 1628
rect 3733 1146 3737 1369
rect 3733 912 3737 1142
rect 3733 684 3737 908
rect 3733 456 3737 680
rect 3733 164 3737 452
rect 3741 1365 3745 1620
rect 3741 1138 3745 1361
rect 3741 904 3745 1134
rect 3741 676 3745 900
rect 3741 448 3745 672
rect 3741 156 3745 444
use 8XOR2  8XOR2_0
timestamp 1746041965
transform 1 0 -112 0 1 972
box 112 -136 910 98
use 8bitADDSUB  8bitADDSUB_0
timestamp 1746041965
transform 1 0 0 0 1 1663
box 0 -138 2337 133
use 8bitAND2  8bitAND2_0
timestamp 1746041965
transform 1 0 5 0 1 1433
box -5 -135 538 92
use 8bitNOR2  8bitNOR2_0
timestamp 1746041965
transform 1 0 0 0 1 736
box 0 -128 446 100
use 8bitOR2  8bitOR2_0
timestamp 1746041965
transform 1 0 0 0 1 1202
box 0 -132 574 96
use BARREL_SHIFT  BARREL_SHIFT_0
timestamp 1746489366
transform 1 0 81 0 1 480
box -81 -164 3602 128
use Comparator8  Comparator8_0
timestamp 1746041965
transform 1 0 4 0 1 48
box -4 -48 2390 268
use Decoder_2x4  Decoder_2x4_0
timestamp 1746041965
transform 1 0 -252 0 1 1433
box -64 -44 125 91
use INV  INV_0
timestamp 1741159900
transform 1 0 -181 0 1 516
box -4 0 20 91
use NAND3  NAND3_0
timestamp 1741221395
transform 1 0 -160 0 1 224
box -5 0 38 91
use NAND3  NAND3_1
timestamp 1741221395
transform 1 0 -165 0 1 516
box -5 0 38 91
use OR2  OR2_0
timestamp 1740126367
transform 1 0 -40 0 1 1700
box -4 0 45 92
use XNOR2  XNOR2_0
timestamp 1746041965
transform 1 0 -404 0 1 1433
box 0 0 96 94
<< labels >>
rlabel metal1 -415 1647 -415 1647 3 A0
rlabel metal1 -415 1639 -415 1639 3 A1
rlabel metal1 -415 1631 -415 1631 3 A2
rlabel metal1 -415 1623 -415 1623 3 A3
rlabel metal1 -415 1615 -415 1615 3 A4
rlabel metal1 -415 1607 -415 1607 3 A5
rlabel metal1 -415 1599 -415 1599 3 A6
rlabel metal1 -415 1591 -415 1591 3 A7
rlabel metal1 -415 1583 -415 1583 3 B0
rlabel metal1 -415 1575 -415 1575 3 B1
rlabel metal1 -415 1567 -415 1567 3 B2
rlabel metal1 -415 1559 -415 1559 3 B3
rlabel metal1 -415 1551 -415 1551 3 B4
rlabel metal1 -415 1543 -415 1543 3 B5
rlabel metal1 -415 1535 -415 1535 3 B6
rlabel metal1 -415 1527 -415 1527 3 B7
rlabel metal1 3743 1678 3743 1678 7 Y0
rlabel metal1 3742 1670 3742 1670 7 Y1
rlabel metal1 3742 1662 3742 1662 7 Y2
rlabel metal1 3741 1654 3741 1654 7 Y3
rlabel metal1 3742 1646 3742 1646 7 Y4
rlabel metal1 3742 1638 3742 1638 7 Y5
rlabel metal1 3742 1630 3742 1630 7 Y6
rlabel m2contact 3743 1622 3743 1622 7 Y7
rlabel metal1 -411 1694 -411 1694 3 func0
rlabel metal1 -411 1686 -411 1686 3 func1
rlabel metal1 -411 1678 -411 1678 3 func2
rlabel metal1 -411 1711 -411 1711 1 VDD
rlabel metal1 -411 1702 -411 1702 1 VSS
rlabel metal1 -414 406 -414 406 1 RorL
rlabel metal1 -414 494 -414 494 1 Sign
rlabel metal1 3743 1686 3743 1686 7 Overflow
rlabel metal2 -4 1672 -4 1672 1 enb0
rlabel metal1 5 1427 5 1427 1 enb1
rlabel metal1 3 1200 3 1200 1 enb2
rlabel metal1 4 970 4 970 1 enb3
rlabel metal1 -4 738 -4 738 1 enb4
rlabel metal1 -4 318 -4 318 1 enb5
rlabel metal1 -10 10 -10 10 1 enb6
rlabel metal1 639 1671 639 1671 1 Cin
rlabel metal1 638 1678 638 1678 1 Bin
rlabel polysilicon 729 1743 729 1743 1 Sbout
rlabel metal1 3477 462 3477 462 1 output2
rlabel metal1 3477 422 3477 422 1 output7
rlabel metal1 3477 430 3477 430 1 output6
rlabel metal1 3477 438 3477 438 1 output5
rlabel metal1 3477 446 3477 446 1 output4
rlabel metal1 3477 454 3477 454 1 output3
rlabel metal1 3477 470 3477 470 1 output1
rlabel metal1 3477 478 3477 478 1 output0
<< end >>
