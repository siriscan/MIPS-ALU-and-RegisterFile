magic
tech scmos
timestamp 1742681920
<< metal1 >>
rect -54 84 -42 88
rect -54 0 -42 4
rect -46 -8 32 -4
rect 36 -8 73 -4
rect 77 -8 114 -4
rect 118 -8 155 -4
rect 159 -8 196 -4
rect 200 -8 237 -4
rect 241 -8 278 -4
rect 282 -8 319 -4
rect -38 -16 48 -12
rect 52 -16 130 -12
rect 134 -16 212 -12
rect 216 -16 294 -12
rect -30 -24 7 -20
rect 11 -24 89 -20
rect 93 -24 171 -20
rect 175 -24 253 -20
rect -22 -32 98 -28
rect 102 -32 139 -28
rect 143 -32 262 -28
rect 266 -32 303 -28
rect -14 -40 16 -36
rect 20 -40 57 -36
rect 61 -40 180 -36
rect 184 -40 221 -36
rect -6 -48 188 -44
rect 192 -48 229 -44
rect 233 -48 270 -44
rect 274 -48 311 -44
rect 2 -56 24 -52
rect 28 -56 65 -52
rect 69 -56 106 -52
rect 110 -56 147 -52
<< m2contact >>
rect 32 55 36 59
rect 73 55 77 59
rect 114 55 118 59
rect 155 55 159 59
rect 196 55 200 59
rect 237 55 241 59
rect 278 55 282 59
rect 319 55 323 59
rect -58 44 -54 48
rect 24 44 28 48
rect 65 44 69 48
rect 106 44 110 48
rect 147 44 151 48
rect 188 44 192 48
rect 229 44 233 48
rect 270 44 274 48
rect 311 44 315 48
rect -42 36 -38 40
rect -26 36 -22 40
rect -10 36 -6 40
rect 16 32 20 36
rect 57 32 61 36
rect 98 32 102 36
rect 139 32 143 36
rect 180 32 184 36
rect 221 32 225 36
rect 262 32 266 36
rect 303 32 307 36
rect 7 20 11 24
rect 48 20 52 24
rect 89 20 93 24
rect 130 20 134 24
rect 171 20 175 24
rect 212 20 216 24
rect 253 20 257 24
rect 294 20 298 24
rect -50 12 -46 16
rect -34 12 -30 16
rect -18 12 -14 16
rect -2 12 2 16
rect 39 12 43 16
rect 80 12 84 16
rect 121 12 125 16
rect 162 12 166 16
rect 203 12 207 16
rect 244 12 248 16
rect 285 12 289 16
rect 326 12 330 16
rect -50 -8 -46 -4
rect 32 -8 36 -4
rect 73 -8 77 -4
rect 114 -8 118 -4
rect 155 -8 159 -4
rect 196 -8 200 -4
rect 237 -8 241 -4
rect 278 -8 282 -4
rect 319 -8 323 -4
rect -42 -16 -38 -12
rect 48 -16 52 -12
rect 130 -16 134 -12
rect 212 -16 216 -12
rect 294 -16 298 -12
rect -34 -24 -30 -20
rect 7 -24 11 -20
rect 89 -24 93 -20
rect 171 -24 175 -20
rect 253 -24 257 -20
rect -26 -32 -22 -28
rect 98 -32 102 -28
rect 139 -32 143 -28
rect 262 -32 266 -28
rect 303 -32 307 -28
rect -18 -40 -14 -36
rect 16 -40 20 -36
rect 57 -40 61 -36
rect 180 -40 184 -36
rect 221 -40 225 -36
rect -10 -48 -6 -44
rect 188 -48 192 -44
rect 229 -48 233 -44
rect 270 -48 274 -44
rect 311 -48 315 -44
rect -2 -56 2 -52
rect 24 -56 28 -52
rect 65 -56 69 -52
rect 106 -56 110 -52
rect 147 -56 151 -52
<< metal2 >>
rect -58 -8 -54 44
rect -50 -4 -46 12
rect -42 -12 -38 36
rect -34 -20 -30 12
rect -26 -28 -22 36
rect -18 -36 -14 12
rect -10 -44 -6 36
rect -2 -52 2 12
rect 7 -20 11 20
rect 16 -36 20 32
rect 24 -52 28 44
rect 32 -4 36 55
rect 39 -64 43 12
rect 48 -12 52 20
rect 57 -36 61 32
rect 65 -52 69 44
rect 73 -4 77 55
rect 80 -64 84 12
rect 89 -20 93 20
rect 98 -28 102 32
rect 106 -52 110 44
rect 114 -4 118 55
rect 121 -64 125 12
rect 130 -12 134 20
rect 139 -28 143 32
rect 147 -52 151 44
rect 155 -4 159 55
rect 162 -64 166 12
rect 171 -20 175 20
rect 180 -36 184 32
rect 188 -44 192 44
rect 196 -4 200 55
rect 203 -64 207 12
rect 212 -12 216 20
rect 221 -36 225 32
rect 229 -44 233 44
rect 237 -4 241 55
rect 244 -64 248 12
rect 253 -20 257 20
rect 262 -28 266 32
rect 270 -44 274 44
rect 278 -4 282 55
rect 285 -64 289 12
rect 294 -12 298 20
rect 303 -28 307 32
rect 311 -44 315 44
rect 319 -4 323 55
rect 326 -64 330 12
use INV  INV_0
timestamp 1741159900
transform 1 0 -60 0 1 0
box -4 0 20 91
use INV  INV_1
timestamp 1741159900
transform 1 0 -44 0 1 0
box -4 0 20 91
use INV  INV_2
timestamp 1741159900
transform 1 0 -28 0 1 0
box -4 0 20 91
use INV  INV_3
timestamp 1741159900
transform 1 0 -12 0 1 0
box -4 0 20 91
use NAND4  NAND4_0
timestamp 1741157784
transform 1 0 4 0 1 0
box -4 0 45 95
use NAND4  NAND4_1
timestamp 1741157784
transform 1 0 45 0 1 0
box -4 0 45 95
use NAND4  NAND4_2
timestamp 1741157784
transform 1 0 86 0 1 0
box -4 0 45 95
use NAND4  NAND4_3
timestamp 1741157784
transform 1 0 127 0 1 0
box -4 0 45 95
use NAND4  NAND4_4
timestamp 1741157784
transform 1 0 168 0 1 0
box -4 0 45 95
use NAND4  NAND4_5
timestamp 1741157784
transform 1 0 209 0 1 0
box -4 0 45 95
use NAND4  NAND4_6
timestamp 1741157784
transform 1 0 250 0 1 0
box -4 0 45 95
use NAND4  NAND4_7
timestamp 1741157784
transform 1 0 291 0 1 0
box -4 0 45 95
<< labels >>
rlabel metal2 -56 -6 -56 -6 1 EN
rlabel metal1 -36 -14 -36 -14 1 S0
rlabel metal1 -20 -30 -20 -30 1 S1
rlabel metal1 -4 -46 -4 -46 1 S2
rlabel metal2 41 -62 41 -62 1 A0
rlabel metal2 82 -62 82 -62 1 A1
rlabel metal2 123 -62 123 -62 1 A2
rlabel metal2 164 -62 164 -62 1 A3
rlabel metal2 205 -62 205 -62 1 A4
rlabel metal2 246 -62 246 -62 1 A5
rlabel metal2 287 -62 287 -62 1 A6
rlabel metal2 328 -62 328 -62 1 A7
rlabel metal1 -52 2 -52 2 1 VSS
rlabel metal1 -49 86 -49 86 1 VDD
<< end >>
