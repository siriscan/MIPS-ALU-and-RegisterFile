magic
tech scmos
timestamp 1746819933
<< nwell >>
rect 3347 2608 3362 2616
rect 3398 2608 3413 2616
rect 3449 2608 3464 2616
rect 3501 2608 3516 2616
rect 4457 2555 4481 2559
rect 4547 2551 4557 2559
rect 4575 2551 4606 2559
rect 5576 2551 5613 2559
rect 5625 2551 5638 2559
rect 5649 2551 5662 2559
rect 5688 2551 5701 2559
rect 5715 2551 5737 2555
rect 4409 2284 4434 2292
rect 4450 2284 4475 2292
rect 4491 2284 4516 2292
rect 4541 2284 4545 2288
rect 4569 2284 4588 2292
rect 3348 2268 3363 2276
rect 3398 2268 3413 2276
rect 3450 2268 3465 2276
rect 4456 2057 4486 2065
rect 4515 2057 4519 2061
rect 3349 1928 3364 1936
rect 3399 1928 3414 1936
rect 3450 1928 3465 1936
rect 3501 1928 3516 1936
rect 4396 1827 4407 1835
rect 4439 1827 4450 1835
rect 4464 1827 4482 1835
rect 4511 1827 4523 1835
rect 4536 1827 4556 1835
rect 3348 1588 3363 1596
rect 3399 1588 3414 1596
rect 3451 1588 3466 1596
rect 3502 1588 3517 1596
rect 4394 1595 4409 1603
rect 4419 1595 4434 1603
rect 4447 1595 4460 1603
rect 4432 1367 4471 1371
rect 4501 1367 4555 1371
rect 4570 1367 4624 1371
rect 4639 1367 4670 1371
rect 5641 1367 5691 1371
rect 5709 1367 5759 1371
rect 5780 1367 5830 1371
rect 3347 1248 3362 1256
rect 3399 1248 3414 1256
rect 3451 1248 3466 1256
rect 3500 1248 3515 1256
rect 4431 1075 4442 1079
rect 4457 1075 4483 1079
rect 4496 1075 4515 1079
rect 4533 1075 4538 1079
rect 4567 1075 4579 1079
rect 4592 1075 4618 1079
rect 4631 1075 4652 1079
rect 4663 1075 4672 1083
rect 5649 1075 5669 1083
rect 5681 1075 5694 1079
rect 5786 1075 5805 1083
rect 5818 1075 5837 1083
rect 3348 908 3363 916
rect 3400 908 3415 916
rect 3450 908 3465 916
rect 3502 908 3517 916
rect 4535 652 4609 656
rect 3347 572 3362 576
rect 3399 568 3414 576
rect 3449 568 3464 576
rect 3501 568 3516 576
rect 1252 236 1256 240
<< metal1 >>
rect 246 2681 7951 2685
rect 310 2673 7959 2677
rect 374 2665 7967 2669
rect 438 2657 7975 2661
rect 502 2649 7983 2653
rect 566 2641 7991 2645
rect 630 2633 7999 2637
rect 694 2625 8007 2629
rect 0 2608 2 2612
rect 215 2608 237 2612
rect 3700 2608 3899 2612
rect 178 2524 183 2528
rect 3709 2524 3879 2528
rect 2 2516 6 2520
rect 2 2500 6 2504
rect 2 2476 6 2480
rect 2 2468 6 2472
rect 2 2460 6 2464
rect 2 2452 6 2456
rect 8011 2451 8015 2455
rect 2 2444 6 2448
rect 8011 2443 8015 2447
rect 2 2436 6 2440
rect 8011 2435 8015 2439
rect 2 2428 6 2432
rect 8011 2427 8015 2431
rect 2 2420 6 2424
rect 8011 2419 8015 2423
rect 3706 2412 3711 2416
rect 3729 2412 3849 2416
rect 3854 2412 3858 2416
rect 8011 2411 8015 2415
rect 3706 2404 3711 2408
rect 3737 2404 3849 2408
rect 3854 2404 3858 2408
rect 8011 2403 8015 2407
rect 3706 2396 3711 2400
rect 3745 2396 3849 2400
rect 3854 2396 3858 2400
rect 8011 2395 8015 2399
rect 3706 2388 3711 2392
rect 3753 2388 3849 2392
rect 3854 2388 3858 2392
rect 8011 2387 8015 2391
rect 3706 2380 3711 2384
rect 3761 2380 3849 2384
rect 3854 2380 3858 2384
rect 3706 2372 3711 2376
rect 3769 2372 3849 2376
rect 3854 2372 3858 2376
rect 3706 2364 3711 2368
rect 3777 2364 3849 2368
rect 3854 2364 3858 2368
rect 3706 2356 3711 2360
rect 3785 2356 3849 2360
rect 3854 2356 3858 2360
rect 3854 2348 3858 2352
rect 3854 2340 3858 2344
rect 3854 2332 3858 2336
rect 3854 2324 3858 2328
rect 3854 2316 3858 2320
rect 3854 2308 3858 2312
rect 3854 2300 3858 2304
rect 3854 2292 3858 2296
rect 12 2176 26 2180
rect 12 2168 26 2172
rect 12 2152 26 2156
rect 12 2136 26 2140
rect 3709 2072 3713 2076
rect 3709 2064 3713 2068
rect 3709 2056 3713 2060
rect 3709 2048 3713 2052
rect 3709 2040 3713 2044
rect 3709 2032 3713 2036
rect 3709 2024 3713 2028
rect 3709 2016 3713 2020
rect 615 1949 617 1953
rect 12 1933 26 1937
rect 12 1917 26 1921
rect 12 1901 26 1905
rect 5058 1743 5062 1747
rect 3709 1732 3713 1736
rect 3709 1724 3713 1728
rect 3709 1716 3713 1720
rect 3709 1708 3713 1712
rect 3709 1700 3713 1704
rect 3709 1692 3713 1696
rect 11 1685 22 1689
rect 3709 1684 3713 1688
rect 3709 1676 3713 1680
rect 11 1669 22 1673
rect 11 1653 22 1657
rect 3708 1392 3712 1396
rect 3708 1384 3712 1388
rect 3708 1376 3712 1380
rect 3708 1368 3712 1372
rect 3708 1360 3712 1364
rect 3708 1352 3712 1356
rect 3708 1344 3712 1348
rect 3708 1336 3712 1340
rect 3857 1067 3895 1071
rect 3710 1052 3714 1056
rect 3710 1044 3714 1048
rect 3710 1036 3714 1040
rect 3710 1028 3714 1032
rect 3710 1020 3714 1024
rect 3710 1012 3714 1016
rect 3710 1004 3714 1008
rect 3710 996 3714 1000
rect 6226 987 6233 991
rect 3709 824 3886 828
rect 3709 712 3713 716
rect 3709 704 3713 708
rect 3709 696 3713 700
rect 3709 688 3713 692
rect 3709 680 3713 684
rect 3709 672 3713 676
rect 3709 664 3713 668
rect 3709 656 3713 660
rect 4611 603 8010 607
rect 3890 568 3893 572
rect 3729 560 3893 564
rect 3737 552 3893 556
rect 3745 544 3893 548
rect 3753 536 3893 540
rect 3761 528 3893 532
rect 3769 520 3893 524
rect 3777 512 3893 516
rect 3785 504 3893 508
rect 3793 496 3893 500
rect 3801 488 3893 492
rect 3809 480 3893 484
rect 3817 472 3893 476
rect 3825 464 3893 468
rect 3833 456 3893 460
rect 3841 448 3894 452
rect 3849 440 3894 444
rect 3707 372 3711 376
rect 3707 364 3711 368
rect 3707 356 3711 360
rect 3707 348 3711 352
rect 3707 340 3711 344
rect 3707 332 3711 336
rect 3707 324 3711 328
rect 3707 316 3711 320
rect 613 136 642 140
<< m2contact >>
rect 242 2681 246 2685
rect 7951 2681 7955 2685
rect 306 2673 310 2677
rect 7959 2673 7963 2677
rect 370 2665 374 2669
rect 7967 2665 7971 2669
rect 434 2657 438 2661
rect 7975 2657 7979 2661
rect 498 2649 502 2653
rect 7983 2649 7987 2653
rect 562 2641 566 2645
rect 7991 2641 7995 2645
rect 626 2633 630 2637
rect 7999 2633 8003 2637
rect 690 2625 694 2629
rect 8007 2625 8011 2629
rect 2 2608 215 2612
rect 249 2608 278 2612
rect 1143 2608 1191 2612
rect 1209 2608 1252 2612
rect 1271 2608 1324 2612
rect 2211 2608 2247 2612
rect 2268 2608 2272 2612
rect 2416 2608 2420 2612
rect 3297 2608 3312 2612
rect 3347 2608 3362 2612
rect 3398 2608 3413 2612
rect 3449 2608 3464 2612
rect 3483 2608 3487 2612
rect 3501 2608 3516 2612
rect 3899 2608 3903 2612
rect 4397 2551 4405 2555
rect 4433 2551 4444 2555
rect 4457 2551 4481 2555
rect 4531 2551 4535 2555
rect 4547 2551 4557 2555
rect 4575 2551 4606 2555
rect 5576 2551 5613 2555
rect 5625 2551 5638 2555
rect 5649 2551 5662 2555
rect 5688 2551 5701 2555
rect 5715 2551 5737 2555
rect 5825 2551 5846 2555
rect 611 2524 615 2528
rect 738 2524 800 2528
rect 1746 2524 1758 2528
rect 1778 2524 1790 2528
rect 1846 2524 1850 2528
rect 2796 2524 2800 2528
rect 2871 2524 2886 2528
rect 2922 2524 2937 2528
rect 3879 2524 3883 2528
rect 3899 2476 3903 2480
rect 3879 2467 3883 2471
rect 3949 2467 4097 2471
rect 5051 2467 5067 2471
rect 5224 2467 5234 2471
rect 6225 2467 6238 2471
rect 6300 2467 6319 2471
rect 6356 2467 6367 2471
rect 3912 2459 3916 2463
rect 3920 2451 3924 2455
rect 3928 2443 3932 2447
rect 3725 2412 3729 2416
rect 3733 2404 3737 2408
rect 3741 2396 3745 2400
rect 3749 2388 3753 2392
rect 3757 2380 3761 2384
rect 3765 2372 3769 2376
rect 3773 2364 3777 2368
rect 3781 2356 3785 2360
rect 4409 2284 4434 2288
rect 4450 2284 4475 2288
rect 4491 2284 4516 2288
rect 4530 2284 4555 2288
rect 4569 2284 4588 2288
rect 4602 2284 4668 2288
rect 2 2268 187 2272
rect 200 2268 206 2272
rect 215 2268 221 2272
rect 231 2268 237 2272
rect 247 2268 262 2272
rect 271 2268 279 2272
rect 1144 2268 1192 2272
rect 1206 2268 1254 2272
rect 1272 2268 1326 2272
rect 2211 2268 2246 2272
rect 2416 2268 2420 2272
rect 3297 2268 3312 2272
rect 3348 2268 3363 2272
rect 3398 2268 3413 2272
rect 3450 2268 3465 2272
rect 3484 2268 3488 2272
rect 3892 2200 3911 2204
rect 795 2184 802 2188
rect 1746 2184 1758 2188
rect 1778 2184 1790 2188
rect 1847 2184 1851 2188
rect 2797 2184 2801 2188
rect 2869 2184 2884 2188
rect 2921 2184 2936 2188
rect 4413 2057 4443 2061
rect 4456 2057 4486 2061
rect 4501 2057 4531 2061
rect 4589 2057 4619 2061
rect 4 2033 217 2037
rect 3944 1973 3967 1977
rect 3982 1973 4052 1977
rect 617 1949 621 1953
rect 1143 1928 1191 1932
rect 1207 1928 1255 1932
rect 1271 1928 1326 1932
rect 2211 1928 2246 1932
rect 2416 1928 2420 1932
rect 3297 1928 3312 1932
rect 3349 1928 3364 1932
rect 3399 1928 3414 1932
rect 3450 1928 3465 1932
rect 3483 1928 3487 1932
rect 3501 1928 3516 1932
rect 576 1844 604 1848
rect 697 1844 712 1848
rect 1746 1844 1758 1848
rect 1778 1844 1790 1848
rect 1848 1844 1852 1848
rect 2796 1844 2800 1848
rect 2869 1844 2884 1848
rect 2921 1844 2936 1848
rect 4396 1827 4407 1831
rect 4439 1827 4450 1831
rect 4464 1827 4482 1831
rect 4511 1827 4523 1831
rect 4536 1827 4556 1831
rect 4609 1827 4627 1831
rect 185 1785 195 1789
rect 225 1785 235 1789
rect 267 1785 277 1789
rect 3943 1743 3966 1747
rect 3980 1743 4087 1747
rect 5062 1743 5066 1747
rect 4394 1595 4409 1599
rect 4419 1595 4434 1599
rect 4447 1595 4460 1599
rect 4477 1595 4490 1599
rect 4506 1595 4510 1599
rect 4 1588 219 1592
rect 1144 1588 1191 1592
rect 1207 1588 1255 1592
rect 1271 1588 1326 1592
rect 2212 1588 2247 1592
rect 2417 1588 2421 1592
rect 3297 1588 3312 1592
rect 3348 1588 3363 1592
rect 3399 1588 3414 1592
rect 3451 1588 3466 1592
rect 3482 1588 3486 1592
rect 3502 1588 3517 1592
rect 3983 1511 4105 1515
rect 578 1504 604 1508
rect 618 1504 636 1508
rect 698 1504 723 1508
rect 1747 1504 1759 1508
rect 1778 1504 1790 1508
rect 1848 1504 1852 1508
rect 2797 1504 2801 1508
rect 2870 1504 2885 1508
rect 2920 1504 2935 1508
rect 4395 1367 4418 1371
rect 4432 1367 4471 1371
rect 4501 1367 4555 1371
rect 4570 1367 4624 1371
rect 4639 1367 4670 1371
rect 5575 1367 5624 1371
rect 5641 1367 5691 1371
rect 5709 1367 5759 1371
rect 5780 1367 5830 1371
rect 6744 1367 6763 1371
rect 6780 1367 6834 1371
rect 6849 1367 6903 1371
rect 6919 1367 6973 1371
rect 6987 1367 7009 1371
rect 3981 1283 4080 1287
rect 5051 1283 5062 1287
rect 5121 1283 5132 1287
rect 5189 1283 5200 1287
rect 5259 1283 5270 1287
rect 6191 1283 6202 1287
rect 6262 1283 6273 1287
rect 6329 1283 6340 1287
rect 6399 1283 6410 1287
rect 7331 1283 7342 1287
rect 7401 1283 7412 1287
rect 7469 1283 7480 1287
rect 7538 1283 7549 1287
rect 3876 1259 3880 1263
rect 7 1248 259 1252
rect 1143 1248 1192 1252
rect 1207 1248 1253 1252
rect 1270 1248 1328 1252
rect 2211 1248 2246 1252
rect 2416 1248 2420 1252
rect 3297 1248 3312 1252
rect 3347 1248 3362 1252
rect 3399 1248 3414 1252
rect 3451 1248 3466 1252
rect 3483 1248 3487 1252
rect 3500 1248 3515 1252
rect 3895 1171 3899 1175
rect 577 1164 600 1168
rect 619 1164 649 1168
rect 698 1164 727 1168
rect 1747 1164 1759 1168
rect 1778 1164 1790 1168
rect 1848 1164 1852 1168
rect 2797 1164 2801 1168
rect 2870 1164 2885 1168
rect 2922 1164 2937 1168
rect 4079 1075 4083 1079
rect 4431 1075 4442 1079
rect 4457 1075 4483 1079
rect 4496 1075 4515 1079
rect 4529 1075 4538 1079
rect 4567 1075 4579 1079
rect 4592 1075 4618 1079
rect 4631 1075 4652 1079
rect 4663 1075 4672 1079
rect 5585 1075 5598 1079
rect 5611 1075 5636 1079
rect 5649 1075 5669 1079
rect 5681 1075 5694 1079
rect 5745 1075 5771 1079
rect 5786 1075 5805 1079
rect 5818 1075 5837 1079
rect 3853 1067 3857 1071
rect 3895 1067 3899 1071
rect 3945 991 4075 995
rect 5034 991 5044 995
rect 5074 991 5090 995
rect 5113 991 5129 995
rect 5152 991 5168 995
rect 6138 991 6149 995
rect 6171 991 6182 995
rect 6226 991 6233 995
rect 6268 991 6272 995
rect 7 908 274 912
rect 1141 908 1191 912
rect 1206 908 1256 912
rect 1269 908 1328 912
rect 2212 908 2247 912
rect 2416 908 2420 912
rect 3296 908 3311 912
rect 3348 908 3363 912
rect 3400 908 3415 912
rect 3450 908 3465 912
rect 3483 908 3487 912
rect 3502 908 3517 912
rect 576 824 604 828
rect 618 824 665 828
rect 699 824 724 828
rect 1746 824 1758 828
rect 1778 824 1790 828
rect 1848 824 1852 828
rect 2797 824 2801 828
rect 2870 824 2885 828
rect 2921 824 2936 828
rect 3886 824 3890 828
rect 4079 652 4083 656
rect 4394 652 4407 656
rect 4418 652 4446 656
rect 4473 652 4487 656
rect 4499 652 4521 656
rect 4535 652 4609 656
rect 6 568 278 572
rect 1142 568 1191 572
rect 1206 568 1255 572
rect 1272 568 1321 572
rect 2212 568 2247 572
rect 2415 568 2419 572
rect 3297 568 3312 572
rect 3347 568 3362 572
rect 3399 568 3414 572
rect 3449 568 3464 572
rect 3483 568 3487 572
rect 3501 568 3516 572
rect 3886 568 3890 572
rect 3921 568 3936 572
rect 3997 568 4012 572
rect 4042 568 4046 572
rect 4078 568 4093 572
rect 3725 560 3729 564
rect 3733 552 3737 556
rect 3741 544 3745 548
rect 3749 536 3753 540
rect 3757 528 3761 532
rect 3765 520 3769 524
rect 3773 512 3777 516
rect 3781 504 3785 508
rect 3789 496 3793 500
rect 3797 488 3801 492
rect 575 484 603 488
rect 617 484 681 488
rect 698 484 726 488
rect 1746 484 1758 488
rect 1777 484 1789 488
rect 1848 484 1852 488
rect 2797 484 2801 488
rect 2870 484 2885 488
rect 2922 484 2937 488
rect 3805 480 3809 484
rect 3813 472 3817 476
rect 3821 464 3825 468
rect 3829 456 3833 460
rect 3837 448 3841 452
rect 3845 440 3849 444
rect 5 236 277 240
rect 1165 236 1180 240
rect 1243 236 1254 240
rect 1268 236 1283 240
rect 569 152 604 156
rect 617 152 634 156
<< metal2 >>
rect 242 2619 246 2681
rect 306 2620 310 2673
rect 370 2619 374 2665
rect 434 2618 438 2657
rect 498 2619 502 2649
rect 562 2620 566 2641
rect 626 2620 630 2633
rect 690 2617 694 2625
rect 3879 2471 3883 2524
rect 3899 2480 3903 2608
rect 3912 2463 3916 2700
rect 3920 2455 3924 2700
rect 3928 2447 3932 2700
rect 7951 2426 7955 2681
rect 7959 2426 7963 2673
rect 7967 2426 7971 2665
rect 7975 2421 7979 2657
rect 3725 2356 3729 2412
rect 3733 2408 3737 2416
rect 3733 2356 3737 2404
rect 3741 2400 3745 2416
rect 3741 2356 3745 2396
rect 3749 2392 3753 2416
rect 3749 2356 3753 2388
rect 3757 2384 3761 2416
rect 3757 2356 3761 2380
rect 3765 2376 3769 2416
rect 3765 2356 3769 2372
rect 3773 2368 3777 2416
rect 3773 2356 3777 2364
rect 3781 2360 3785 2416
rect 7983 2394 7987 2649
rect 7991 2399 7995 2641
rect 7999 2392 8003 2633
rect 8007 2391 8011 2625
rect 3725 440 3729 560
rect 3733 556 3737 564
rect 3733 440 3737 552
rect 3741 548 3745 564
rect 3741 440 3745 544
rect 3749 540 3753 564
rect 3749 440 3753 536
rect 3757 532 3761 564
rect 3757 440 3761 528
rect 3765 524 3769 564
rect 3765 440 3769 520
rect 3773 516 3777 564
rect 3773 440 3777 512
rect 3781 508 3785 564
rect 3781 440 3785 504
rect 3789 500 3793 564
rect 3789 440 3793 496
rect 3797 492 3801 564
rect 3797 440 3801 488
rect 3805 484 3809 564
rect 3805 440 3809 480
rect 3813 476 3817 564
rect 3813 440 3817 472
rect 3821 468 3825 564
rect 3821 440 3825 464
rect 3829 460 3833 564
rect 3829 440 3833 456
rect 3837 452 3841 564
rect 3837 440 3841 448
rect 3845 444 3849 564
rect 3853 -12 3857 1067
rect 3876 -12 3880 1259
rect 3895 1071 3899 1171
rect 3886 572 3890 824
rect 4079 656 4083 1075
<< m3contact >>
rect 2 2612 215 2616
rect 249 2612 278 2616
rect 1143 2612 1191 2616
rect 1209 2612 1252 2616
rect 1271 2612 1324 2616
rect 2211 2612 2247 2616
rect 2416 2612 2420 2616
rect 3297 2612 3312 2616
rect 3347 2612 3362 2616
rect 3398 2612 3413 2616
rect 3449 2612 3464 2616
rect 3501 2612 3516 2616
rect 3483 2604 3487 2608
rect 738 2528 800 2532
rect 1846 2528 1850 2532
rect 615 2524 619 2528
rect 1746 2520 1758 2524
rect 2796 2528 2800 2532
rect 1778 2520 1790 2524
rect 2871 2520 2886 2524
rect 2922 2520 2937 2524
rect 4397 2555 4405 2559
rect 4433 2555 4444 2559
rect 4457 2555 4481 2559
rect 4531 2555 4535 2559
rect 4547 2555 4557 2559
rect 4575 2555 4606 2559
rect 5576 2555 5613 2559
rect 5625 2555 5638 2559
rect 5649 2555 5662 2559
rect 5688 2555 5701 2559
rect 5715 2555 5737 2559
rect 5825 2555 5846 2559
rect 3949 2471 4097 2475
rect 5051 2463 5067 2467
rect 5224 2463 5234 2467
rect 6225 2463 6238 2467
rect 6300 2463 6319 2467
rect 6356 2463 6367 2467
rect 4409 2288 4434 2292
rect 4450 2288 4475 2292
rect 4491 2288 4516 2292
rect 4530 2288 4555 2292
rect 4569 2288 4588 2292
rect 4602 2288 4668 2292
rect 2 2272 187 2276
rect 200 2272 206 2276
rect 215 2272 221 2276
rect 231 2272 237 2276
rect 247 2272 262 2276
rect 271 2272 279 2276
rect 1144 2272 1192 2276
rect 1206 2272 1254 2276
rect 1272 2272 1326 2276
rect 2211 2272 2246 2276
rect 2416 2272 2420 2276
rect 3297 2272 3312 2276
rect 3348 2272 3363 2276
rect 3398 2272 3413 2276
rect 3450 2272 3465 2276
rect 3484 2264 3488 2268
rect 3892 2196 3911 2200
rect 795 2188 802 2192
rect 1847 2188 1851 2192
rect 1746 2180 1758 2184
rect 2797 2188 2801 2192
rect 1778 2180 1790 2184
rect 2869 2180 2884 2184
rect 2921 2180 2936 2184
rect 4413 2061 4443 2065
rect 4456 2061 4486 2065
rect 4501 2061 4531 2065
rect 4589 2061 4619 2065
rect 4 2037 217 2041
rect 3944 1977 3967 1981
rect 3982 1977 4052 1981
rect 617 1953 621 1957
rect 1143 1932 1191 1936
rect 1207 1932 1255 1936
rect 1271 1932 1326 1936
rect 2211 1932 2246 1936
rect 2416 1932 2420 1936
rect 3297 1932 3312 1936
rect 3349 1932 3364 1936
rect 3399 1932 3414 1936
rect 3450 1932 3465 1936
rect 3501 1932 3516 1936
rect 3483 1924 3487 1928
rect 576 1848 604 1852
rect 697 1848 712 1852
rect 1848 1848 1852 1852
rect 1746 1840 1758 1844
rect 2796 1848 2800 1852
rect 1778 1840 1790 1844
rect 2869 1840 2884 1844
rect 2921 1840 2936 1844
rect 4396 1831 4407 1835
rect 4439 1831 4450 1835
rect 4464 1831 4482 1835
rect 4511 1831 4523 1835
rect 4536 1831 4556 1835
rect 4609 1831 4627 1835
rect 185 1789 195 1793
rect 225 1789 235 1793
rect 267 1789 277 1793
rect 3943 1747 3966 1751
rect 3980 1747 4087 1751
rect 5062 1739 5066 1743
rect 4394 1599 4409 1603
rect 4 1592 219 1596
rect 1144 1592 1191 1596
rect 1207 1592 1255 1596
rect 1271 1592 1326 1596
rect 2212 1592 2247 1596
rect 2417 1592 2421 1596
rect 3297 1592 3312 1596
rect 3348 1592 3363 1596
rect 3399 1592 3414 1596
rect 3451 1592 3466 1596
rect 3502 1592 3517 1596
rect 4419 1599 4434 1603
rect 4447 1599 4460 1603
rect 4477 1599 4490 1603
rect 4510 1595 4514 1599
rect 3482 1584 3486 1588
rect 3983 1515 4105 1519
rect 578 1508 604 1512
rect 618 1508 636 1512
rect 698 1508 723 1512
rect 1848 1508 1852 1512
rect 1747 1500 1759 1504
rect 2797 1508 2801 1512
rect 1778 1500 1790 1504
rect 2870 1500 2885 1504
rect 2920 1500 2935 1504
rect 4395 1371 4418 1375
rect 4432 1371 4471 1375
rect 4501 1371 4555 1375
rect 4570 1371 4624 1375
rect 4639 1371 4670 1375
rect 5575 1371 5624 1375
rect 5641 1371 5691 1375
rect 5709 1371 5759 1375
rect 5780 1371 5830 1375
rect 6744 1371 6763 1375
rect 6780 1371 6834 1375
rect 6849 1371 6903 1375
rect 6919 1371 6973 1375
rect 6987 1371 7009 1375
rect 3981 1287 4080 1291
rect 5051 1279 5062 1283
rect 5121 1279 5132 1283
rect 5189 1279 5200 1283
rect 5259 1279 5270 1283
rect 6191 1279 6202 1283
rect 6262 1279 6273 1283
rect 6329 1279 6340 1283
rect 6399 1279 6410 1283
rect 7331 1279 7342 1283
rect 7401 1279 7412 1283
rect 7469 1279 7480 1283
rect 7538 1279 7549 1283
rect 7 1252 259 1256
rect 1143 1252 1192 1256
rect 1207 1252 1253 1256
rect 1270 1252 1328 1256
rect 2211 1252 2246 1256
rect 2416 1252 2420 1256
rect 3297 1252 3312 1256
rect 3347 1252 3362 1256
rect 3399 1252 3414 1256
rect 3451 1252 3466 1256
rect 3500 1252 3515 1256
rect 3483 1244 3487 1248
rect 577 1168 600 1172
rect 619 1168 649 1172
rect 698 1168 727 1172
rect 1848 1168 1852 1172
rect 1747 1160 1759 1164
rect 2797 1168 2801 1172
rect 1778 1160 1790 1164
rect 2870 1160 2885 1164
rect 2922 1160 2937 1164
rect 7 912 274 916
rect 1141 912 1191 916
rect 1206 912 1256 916
rect 1269 912 1328 916
rect 2212 912 2247 916
rect 2416 912 2420 916
rect 3296 912 3311 916
rect 3348 912 3363 916
rect 3400 912 3415 916
rect 3450 912 3465 916
rect 3502 912 3517 916
rect 3483 904 3487 908
rect 576 828 604 832
rect 618 828 665 832
rect 699 828 724 832
rect 1848 828 1852 832
rect 1746 820 1758 824
rect 2797 828 2801 832
rect 1778 820 1790 824
rect 2870 820 2885 824
rect 2921 820 2936 824
rect 6 572 278 576
rect 1142 572 1191 576
rect 1206 572 1255 576
rect 1272 572 1321 576
rect 2212 572 2247 576
rect 2415 572 2419 576
rect 3297 572 3312 576
rect 3347 572 3362 576
rect 3399 572 3414 576
rect 3449 572 3464 576
rect 3501 572 3516 576
rect 3483 564 3487 568
rect 575 488 603 492
rect 617 488 681 492
rect 698 488 726 492
rect 1848 488 1852 492
rect 1746 480 1758 484
rect 2797 488 2801 492
rect 1777 480 1789 484
rect 2870 480 2885 484
rect 2922 480 2937 484
rect 5 240 277 244
rect 1165 240 1180 244
rect 1243 240 1254 244
rect 1268 240 1283 244
rect 569 156 604 160
rect 617 156 634 160
rect 4431 1079 4442 1083
rect 4457 1079 4483 1083
rect 4496 1079 4515 1083
rect 4529 1079 4538 1083
rect 4567 1079 4579 1083
rect 4592 1079 4618 1083
rect 4631 1079 4652 1083
rect 4663 1079 4672 1083
rect 5585 1079 5598 1083
rect 5611 1079 5636 1083
rect 5649 1079 5669 1083
rect 5681 1079 5694 1083
rect 5745 1079 5771 1083
rect 5786 1079 5805 1083
rect 5818 1079 5837 1083
rect 3945 995 4075 999
rect 5034 987 5044 991
rect 5074 987 5090 991
rect 5113 987 5129 991
rect 5152 987 5168 991
rect 6138 987 6149 991
rect 6171 987 6182 991
rect 6226 987 6233 991
rect 6268 987 6272 991
rect 4394 656 4407 660
rect 4418 656 4446 660
rect 4473 656 4487 660
rect 4499 656 4521 660
rect 4535 656 4609 660
rect 4042 572 4046 576
rect 3921 564 3936 568
rect 3997 564 4012 568
rect 4078 564 4093 568
<< metal3 >>
rect -10 3141 8178 3326
rect -32 2958 8178 3141
rect -32 2930 8172 2958
rect -32 2926 502 2930
rect 921 2928 8172 2930
rect 921 2927 7188 2928
rect 921 2926 3745 2927
rect 4164 2926 7188 2927
rect 7607 2926 8172 2928
rect 0 2616 282 2926
rect 0 2612 2 2616
rect 215 2612 249 2616
rect 278 2612 282 2616
rect 0 2276 282 2612
rect 0 2272 2 2276
rect 187 2272 200 2276
rect 206 2272 215 2276
rect 221 2272 231 2276
rect 237 2272 247 2276
rect 262 2272 271 2276
rect 279 2272 282 2276
rect 0 2041 282 2272
rect 0 2037 4 2041
rect 217 2037 282 2041
rect 0 1793 282 2037
rect 0 1789 185 1793
rect 195 1789 225 1793
rect 235 1789 267 1793
rect 277 1789 282 1793
rect 0 1596 282 1789
rect 0 1592 4 1596
rect 219 1592 282 1596
rect 0 1256 282 1592
rect 0 1252 7 1256
rect 259 1252 282 1256
rect 0 916 282 1252
rect 0 912 7 916
rect 274 912 282 916
rect 0 576 282 912
rect 0 572 6 576
rect 278 572 282 576
rect 0 244 282 572
rect 0 240 5 244
rect 277 240 282 244
rect 0 148 282 240
rect 566 2532 848 2737
rect 566 2528 738 2532
rect 800 2528 848 2532
rect 566 2524 615 2528
rect 619 2524 848 2528
rect 566 2192 848 2524
rect 566 2188 795 2192
rect 802 2188 848 2192
rect 566 1957 848 2188
rect 566 1953 617 1957
rect 621 1953 848 1957
rect 566 1852 848 1953
rect 566 1848 576 1852
rect 604 1848 697 1852
rect 712 1848 848 1852
rect 566 1512 848 1848
rect 566 1508 578 1512
rect 604 1508 618 1512
rect 636 1508 698 1512
rect 723 1508 848 1512
rect 566 1172 848 1508
rect 566 1168 577 1172
rect 600 1168 619 1172
rect 649 1168 698 1172
rect 727 1168 848 1172
rect 566 832 848 1168
rect 566 828 576 832
rect 604 828 618 832
rect 665 828 699 832
rect 724 828 848 832
rect 566 492 848 828
rect 566 488 575 492
rect 603 488 617 492
rect 681 488 698 492
rect 726 488 848 492
rect 566 160 848 488
rect 566 156 569 160
rect 604 156 617 160
rect 634 156 848 160
rect 566 18 848 156
rect 1129 2616 1411 2926
rect 1129 2612 1143 2616
rect 1191 2612 1209 2616
rect 1252 2612 1271 2616
rect 1324 2612 1411 2616
rect 1129 2276 1411 2612
rect 1129 2272 1144 2276
rect 1192 2272 1206 2276
rect 1254 2272 1272 2276
rect 1326 2272 1411 2276
rect 1129 1936 1411 2272
rect 1129 1932 1143 1936
rect 1191 1932 1207 1936
rect 1255 1932 1271 1936
rect 1326 1932 1411 1936
rect 1129 1596 1411 1932
rect 1129 1592 1144 1596
rect 1191 1592 1207 1596
rect 1255 1592 1271 1596
rect 1326 1592 1411 1596
rect 1129 1256 1411 1592
rect 1129 1252 1143 1256
rect 1192 1252 1207 1256
rect 1253 1252 1270 1256
rect 1328 1252 1411 1256
rect 1129 916 1411 1252
rect 1129 912 1141 916
rect 1191 912 1206 916
rect 1256 912 1269 916
rect 1328 912 1411 916
rect 1129 576 1411 912
rect 1129 572 1142 576
rect 1191 572 1206 576
rect 1255 572 1272 576
rect 1321 572 1411 576
rect 1129 244 1411 572
rect 1129 240 1165 244
rect 1180 240 1243 244
rect 1254 240 1268 244
rect 1283 240 1411 244
rect 1129 142 1411 240
rect 1616 2532 1889 2733
rect 1616 2528 1846 2532
rect 1850 2528 1889 2532
rect 1616 2524 1889 2528
rect 1616 2520 1746 2524
rect 1758 2520 1778 2524
rect 1790 2520 1889 2524
rect 1616 2192 1889 2520
rect 1616 2188 1847 2192
rect 1851 2188 1889 2192
rect 1616 2184 1889 2188
rect 1616 2180 1746 2184
rect 1758 2180 1778 2184
rect 1790 2180 1889 2184
rect 1616 1852 1889 2180
rect 1616 1848 1848 1852
rect 1852 1848 1889 1852
rect 1616 1844 1889 1848
rect 1616 1840 1746 1844
rect 1758 1840 1778 1844
rect 1790 1840 1889 1844
rect 1616 1512 1889 1840
rect 1616 1508 1848 1512
rect 1852 1508 1889 1512
rect 1616 1504 1889 1508
rect 1616 1500 1747 1504
rect 1759 1500 1778 1504
rect 1790 1500 1889 1504
rect 1616 1172 1889 1500
rect 1616 1168 1848 1172
rect 1852 1168 1889 1172
rect 1616 1164 1889 1168
rect 1616 1160 1747 1164
rect 1759 1160 1778 1164
rect 1790 1160 1889 1164
rect 1616 832 1889 1160
rect 1616 828 1848 832
rect 1852 828 1889 832
rect 1616 824 1889 828
rect 1616 820 1746 824
rect 1758 820 1778 824
rect 1790 820 1889 824
rect 1616 492 1889 820
rect 1616 488 1848 492
rect 1852 488 1889 492
rect 1616 484 1889 488
rect 1616 480 1746 484
rect 1758 480 1777 484
rect 1789 480 1889 484
rect 1616 18 1889 480
rect 2173 2616 2455 2926
rect 2173 2612 2211 2616
rect 2247 2612 2416 2616
rect 2420 2612 2455 2616
rect 2173 2276 2455 2612
rect 2173 2272 2211 2276
rect 2246 2272 2416 2276
rect 2420 2272 2455 2276
rect 2173 1936 2455 2272
rect 2173 1932 2211 1936
rect 2246 1932 2416 1936
rect 2420 1932 2455 1936
rect 2173 1596 2455 1932
rect 2173 1592 2212 1596
rect 2247 1592 2417 1596
rect 2421 1592 2455 1596
rect 2173 1256 2455 1592
rect 2173 1252 2211 1256
rect 2246 1252 2416 1256
rect 2420 1252 2455 1256
rect 2173 916 2455 1252
rect 2173 912 2212 916
rect 2247 912 2416 916
rect 2420 912 2455 916
rect 2173 576 2455 912
rect 2173 572 2212 576
rect 2247 572 2415 576
rect 2419 572 2455 576
rect 2173 139 2455 572
rect 2736 2532 3018 2733
rect 2736 2528 2796 2532
rect 2800 2528 3018 2532
rect 2736 2524 3018 2528
rect 2736 2520 2871 2524
rect 2886 2520 2922 2524
rect 2937 2520 3018 2524
rect 2736 2192 3018 2520
rect 2736 2188 2797 2192
rect 2801 2188 3018 2192
rect 2736 2184 3018 2188
rect 2736 2180 2869 2184
rect 2884 2180 2921 2184
rect 2936 2180 3018 2184
rect 2736 1852 3018 2180
rect 2736 1848 2796 1852
rect 2800 1848 3018 1852
rect 2736 1844 3018 1848
rect 2736 1840 2869 1844
rect 2884 1840 2921 1844
rect 2936 1840 3018 1844
rect 2736 1512 3018 1840
rect 2736 1508 2797 1512
rect 2801 1508 3018 1512
rect 2736 1504 3018 1508
rect 2736 1500 2870 1504
rect 2885 1500 2920 1504
rect 2935 1500 3018 1504
rect 2736 1172 3018 1500
rect 2736 1168 2797 1172
rect 2801 1168 3018 1172
rect 2736 1164 3018 1168
rect 2736 1160 2870 1164
rect 2885 1160 2922 1164
rect 2937 1160 3018 1164
rect 2736 832 3018 1160
rect 2736 828 2797 832
rect 2801 828 3018 832
rect 2736 824 3018 828
rect 2736 820 2870 824
rect 2885 820 2921 824
rect 2936 820 3018 824
rect 2736 492 3018 820
rect 2736 488 2797 492
rect 2801 488 3018 492
rect 2736 484 3018 488
rect 2736 480 2870 484
rect 2885 480 2922 484
rect 2937 480 3018 484
rect 2736 18 3018 480
rect 3272 2616 3545 2926
rect 3272 2612 3297 2616
rect 3312 2612 3347 2616
rect 3362 2612 3398 2616
rect 3413 2612 3449 2616
rect 3464 2612 3501 2616
rect 3516 2612 3545 2616
rect 3272 2608 3545 2612
rect 3272 2604 3483 2608
rect 3487 2604 3545 2608
rect 3272 2276 3545 2604
rect 3272 2272 3297 2276
rect 3312 2272 3348 2276
rect 3363 2272 3398 2276
rect 3413 2272 3450 2276
rect 3465 2272 3545 2276
rect 3272 2268 3545 2272
rect 3272 2264 3484 2268
rect 3488 2264 3545 2268
rect 3272 1936 3545 2264
rect 3272 1932 3297 1936
rect 3312 1932 3349 1936
rect 3364 1932 3399 1936
rect 3414 1932 3450 1936
rect 3465 1932 3501 1936
rect 3516 1932 3545 1936
rect 3272 1928 3545 1932
rect 3272 1924 3483 1928
rect 3487 1924 3545 1928
rect 3272 1596 3545 1924
rect 3272 1592 3297 1596
rect 3312 1592 3348 1596
rect 3363 1592 3399 1596
rect 3414 1592 3451 1596
rect 3466 1592 3502 1596
rect 3517 1592 3545 1596
rect 3272 1588 3545 1592
rect 3272 1584 3482 1588
rect 3486 1584 3545 1588
rect 3272 1256 3545 1584
rect 3272 1252 3297 1256
rect 3312 1252 3347 1256
rect 3362 1252 3399 1256
rect 3414 1252 3451 1256
rect 3466 1252 3500 1256
rect 3515 1252 3545 1256
rect 3272 1248 3545 1252
rect 3272 1244 3483 1248
rect 3487 1244 3545 1248
rect 3272 916 3545 1244
rect 3272 912 3296 916
rect 3311 912 3348 916
rect 3363 912 3400 916
rect 3415 912 3450 916
rect 3465 912 3502 916
rect 3517 912 3545 916
rect 3272 908 3545 912
rect 3272 904 3483 908
rect 3487 904 3545 908
rect 3272 576 3545 904
rect 3272 572 3297 576
rect 3312 572 3347 576
rect 3362 572 3399 576
rect 3414 572 3449 576
rect 3464 572 3501 576
rect 3516 572 3545 576
rect 3272 568 3545 572
rect 3272 564 3483 568
rect 3487 564 3545 568
rect 3272 150 3545 564
rect 3829 2475 4111 2734
rect 3829 2471 3949 2475
rect 4097 2471 4111 2475
rect 3829 2200 4111 2471
rect 3829 2196 3892 2200
rect 3911 2196 4111 2200
rect 3829 1981 4111 2196
rect 3829 1977 3944 1981
rect 3967 1977 3982 1981
rect 4052 1977 4111 1981
rect 3829 1751 4111 1977
rect 3829 1747 3943 1751
rect 3966 1747 3980 1751
rect 4087 1747 4111 1751
rect 3829 1519 4111 1747
rect 3829 1515 3983 1519
rect 4105 1515 4111 1519
rect 3829 1291 4111 1515
rect 3829 1287 3981 1291
rect 4080 1287 4111 1291
rect 3829 999 4111 1287
rect 3829 995 3945 999
rect 4075 995 4111 999
rect 3829 576 4111 995
rect 3829 572 4042 576
rect 4046 572 4111 576
rect 3829 568 4111 572
rect 3829 564 3921 568
rect 3936 564 3997 568
rect 4012 564 4078 568
rect 4093 564 4111 568
rect 3829 18 4111 564
rect 4392 2559 4674 2926
rect 5011 2922 5284 2926
rect 4392 2555 4397 2559
rect 4405 2555 4433 2559
rect 4444 2555 4457 2559
rect 4481 2555 4531 2559
rect 4535 2555 4547 2559
rect 4557 2555 4575 2559
rect 4606 2555 4674 2559
rect 4392 2292 4674 2555
rect 4392 2288 4409 2292
rect 4434 2288 4450 2292
rect 4475 2288 4491 2292
rect 4516 2288 4530 2292
rect 4555 2288 4569 2292
rect 4588 2288 4602 2292
rect 4668 2288 4674 2292
rect 4392 2065 4674 2288
rect 4392 2061 4413 2065
rect 4443 2061 4456 2065
rect 4486 2061 4501 2065
rect 4531 2061 4589 2065
rect 4619 2061 4674 2065
rect 4392 1835 4674 2061
rect 4392 1831 4396 1835
rect 4407 1831 4439 1835
rect 4450 1831 4464 1835
rect 4482 1831 4511 1835
rect 4523 1831 4536 1835
rect 4556 1831 4609 1835
rect 4627 1831 4674 1835
rect 4392 1603 4674 1831
rect 4392 1599 4394 1603
rect 4409 1599 4419 1603
rect 4434 1599 4447 1603
rect 4460 1599 4477 1603
rect 4490 1599 4674 1603
rect 4392 1595 4510 1599
rect 4514 1595 4674 1599
rect 4392 1375 4674 1595
rect 4392 1371 4395 1375
rect 4418 1371 4432 1375
rect 4471 1371 4501 1375
rect 4555 1371 4570 1375
rect 4624 1371 4639 1375
rect 4670 1371 4674 1375
rect 4392 1083 4674 1371
rect 4392 1079 4431 1083
rect 4442 1079 4457 1083
rect 4483 1079 4496 1083
rect 4515 1079 4529 1083
rect 4538 1079 4567 1083
rect 4579 1079 4592 1083
rect 4618 1079 4631 1083
rect 4652 1079 4663 1083
rect 4672 1079 4674 1083
rect 4392 660 4674 1079
rect 4392 656 4394 660
rect 4407 656 4418 660
rect 4446 656 4473 660
rect 4487 656 4499 660
rect 4521 656 4535 660
rect 4609 656 4674 660
rect 4392 141 4674 656
rect 5011 2467 5284 2729
rect 5011 2463 5051 2467
rect 5067 2463 5224 2467
rect 5234 2463 5284 2467
rect 5011 1743 5284 2463
rect 5011 1739 5062 1743
rect 5066 1739 5284 1743
rect 5011 1283 5284 1739
rect 5011 1279 5051 1283
rect 5062 1279 5121 1283
rect 5132 1279 5189 1283
rect 5200 1279 5259 1283
rect 5270 1279 5284 1283
rect 5011 991 5284 1279
rect 5011 987 5034 991
rect 5044 987 5074 991
rect 5090 987 5113 991
rect 5129 987 5152 991
rect 5168 987 5284 991
rect 5011 18 5284 987
rect 5568 2559 5850 2926
rect 6131 2924 6413 2926
rect 5568 2555 5576 2559
rect 5613 2555 5625 2559
rect 5638 2555 5649 2559
rect 5662 2555 5688 2559
rect 5701 2555 5715 2559
rect 5737 2555 5825 2559
rect 5846 2555 5850 2559
rect 5568 1375 5850 2555
rect 5568 1371 5575 1375
rect 5624 1371 5641 1375
rect 5691 1371 5709 1375
rect 5759 1371 5780 1375
rect 5830 1371 5850 1375
rect 5568 1083 5850 1371
rect 5568 1079 5585 1083
rect 5598 1079 5611 1083
rect 5636 1079 5649 1083
rect 5669 1079 5681 1083
rect 5694 1079 5745 1083
rect 5771 1079 5786 1083
rect 5805 1079 5818 1083
rect 5837 1079 5850 1083
rect 5568 141 5850 1079
rect 6131 2467 6413 2731
rect 6131 2463 6225 2467
rect 6238 2463 6300 2467
rect 6319 2463 6356 2467
rect 6367 2463 6413 2467
rect 6131 1283 6413 2463
rect 6131 1279 6191 1283
rect 6202 1279 6262 1283
rect 6273 1279 6329 1283
rect 6340 1279 6399 1283
rect 6410 1279 6413 1283
rect 6131 991 6413 1279
rect 6131 987 6138 991
rect 6149 987 6171 991
rect 6182 987 6226 991
rect 6233 987 6268 991
rect 6272 987 6413 991
rect 6131 18 6413 987
rect 6739 1375 7012 2926
rect 6739 1371 6744 1375
rect 6763 1371 6780 1375
rect 6834 1371 6849 1375
rect 6903 1371 6919 1375
rect 6973 1371 6987 1375
rect 7009 1371 7012 1375
rect 6739 152 7012 1371
rect 7296 1283 7578 2735
rect 7296 1279 7331 1283
rect 7342 1279 7401 1283
rect 7412 1279 7469 1283
rect 7480 1279 7538 1283
rect 7549 1279 7578 1283
rect 7296 33 7578 1279
rect 7859 155 8141 2926
rect 7290 18 7587 33
rect -4 -13 8201 18
rect -6 -420 8201 -13
use ALU  ALU_0
timestamp 1746750801
transform 1 0 4266 0 1 767
box -417 0 3745 1796
use EQUALv2  EQUALv2_0
timestamp 1746688264
transform 1 0 3889 0 1 568
box 0 -128 733 94
use REGISTER_FILEv2  REGISTER_FILEv2_0
timestamp 1746770961
transform 1 0 791 0 1 2276
box -807 -2276 3058 345
<< labels >>
rlabel metal1 180 2526 180 2526 1 VSS
rlabel metal1 3855 2414 3855 2414 3 A0
rlabel metal1 3855 2406 3855 2406 3 A1
rlabel metal1 3855 2398 3855 2398 3 A2
rlabel metal1 3855 2390 3855 2390 3 A3
rlabel metal1 3855 2382 3855 2382 3 A4
rlabel metal1 3855 2374 3855 2374 3 A5
rlabel metal1 3855 2366 3855 2366 3 A6
rlabel metal1 3855 2358 3855 2358 3 A7
rlabel metal1 3855 2350 3855 2350 3 B0
rlabel metal1 3855 2342 3855 2342 3 B1
rlabel metal1 3855 2334 3855 2334 3 B2
rlabel metal1 3855 2326 3855 2326 3 B3
rlabel metal1 3855 2318 3855 2318 3 B4
rlabel metal1 3855 2310 3855 2310 3 B5
rlabel metal1 3855 2302 3855 2302 3 B6
rlabel metal1 3855 2294 3855 2294 3 B7
rlabel metal2 3914 2698 3914 2698 5 func0
rlabel metal2 3922 2698 3922 2698 5 func1
rlabel metal2 3930 2698 3930 2698 5 func2
rlabel metal1 4 2518 4 2518 3 imm_en
rlabel metal1 4 2478 4 2478 1 Imm0
rlabel metal1 4 2470 4 2470 1 Imm1
rlabel metal1 4 2462 4 2462 1 Imm2
rlabel metal1 4 2454 4 2454 1 Imm3
rlabel metal1 4 2446 4 2446 1 Imm4
rlabel metal1 4 2438 4 2438 1 Imm5
rlabel metal1 4 2430 4 2430 1 Imm6
rlabel metal1 4 2422 4 2422 1 Imm7
rlabel space 10 3855 10 3855 5 RorL
rlabel metal2 3878 -10 3878 -10 1 LorA
rlabel metal1 17 2178 17 2178 1 Write_Address3
rlabel metal1 17 2170 17 2170 1 Write_Address0
rlabel metal1 17 2154 17 2154 1 Write_Address1
rlabel metal1 17 2138 17 2138 1 Write_Address2
rlabel metal1 17 1935 17 1935 1 A_Read_Address0
rlabel metal1 17 1919 17 1919 1 A_Read_Address1
rlabel metal1 17 1903 17 1903 1 A_Read_Address2
rlabel metal1 14 1687 14 1687 1 B_Read_Address0
rlabel metal1 14 1671 14 1671 1 B_Read_Address1
rlabel metal1 14 1655 14 1655 1 B_Read_Address2
rlabel metal1 4 2502 4 2502 3 clk
rlabel metal1 3708 2414 3708 2414 1 reg_zero0
rlabel metal1 3708 2406 3708 2406 1 reg_zero1
rlabel metal1 3708 2398 3708 2398 1 reg_zero2
rlabel metal1 3708 2390 3708 2390 1 reg_zero3
rlabel metal1 3708 2382 3708 2382 1 reg_zero4
rlabel metal1 3708 2374 3708 2374 1 reg_zero5
rlabel metal1 3708 2366 3708 2366 1 reg_zero6
rlabel metal1 3708 2358 3708 2358 1 reg_zero7
rlabel metal1 3712 2074 3712 2074 1 reg_one0
rlabel metal1 3712 2066 3712 2066 1 reg_one1
rlabel metal1 3712 2058 3712 2058 1 reg_one2
rlabel metal1 3712 2050 3712 2050 1 reg_one3
rlabel metal1 3712 2042 3712 2042 1 reg_one4
rlabel metal1 3712 2034 3712 2034 1 reg_one5
rlabel metal1 3712 2026 3712 2026 1 reg_one6
rlabel metal1 3712 2018 3712 2018 1 reg_one7
rlabel metal1 3712 1734 3712 1734 1 reg_two0
rlabel metal1 3712 1726 3712 1726 1 reg_two1
rlabel metal1 3712 1718 3712 1718 1 reg_two2
rlabel metal1 3712 1710 3712 1710 1 reg_two3
rlabel metal1 3711 1702 3711 1702 1 reg_two4
rlabel metal1 3712 1694 3712 1694 1 reg_two5
rlabel metal1 3712 1686 3712 1686 1 reg_two6
rlabel metal1 3712 1678 3712 1678 1 reg_two7
rlabel metal1 3711 1394 3711 1394 1 reg_three0
rlabel metal1 3711 1386 3711 1386 1 reg_three1
rlabel metal1 3711 1378 3711 1378 1 reg_three2
rlabel metal1 3711 1370 3711 1370 1 reg_three3
rlabel metal1 3711 1362 3711 1362 1 reg_three4
rlabel metal1 3711 1354 3711 1354 1 reg_three5
rlabel metal1 3711 1346 3711 1346 1 reg_three6
rlabel metal1 3711 1338 3711 1338 1 reg_three7
rlabel metal1 3713 1054 3713 1054 1 reg_four0
rlabel metal1 3713 1046 3713 1046 1 reg_four1
rlabel metal1 3713 1038 3713 1038 1 reg_four2
rlabel metal1 3713 1030 3713 1030 1 reg_four3
rlabel metal1 3713 1022 3713 1022 1 reg_four4
rlabel metal1 3713 1014 3713 1014 1 reg_four5
rlabel metal1 3714 1006 3714 1006 1 reg_four6
rlabel metal1 3714 998 3714 998 1 reg_four7
rlabel metal1 3713 714 3713 714 1 reg_five0
rlabel metal1 3713 706 3713 706 1 reg_five1
rlabel metal1 3712 698 3712 698 1 reg_five2
rlabel metal1 3712 690 3712 690 1 reg_five3
rlabel metal1 3712 682 3712 682 1 reg_five4
rlabel metal1 3712 674 3712 674 1 reg_five5
rlabel metal1 3712 666 3712 666 1 reg_five6
rlabel metal1 3712 658 3712 658 1 reg_five7
rlabel metal1 3710 374 3710 374 1 reg_six0
rlabel metal1 3710 366 3710 366 1 reg_six1
rlabel metal1 3710 358 3710 358 1 reg_six2
rlabel metal1 3710 350 3710 350 1 reg_six3
rlabel metal1 3710 342 3710 342 1 reg_six4
rlabel metal1 3710 334 3710 334 1 reg_six5
rlabel metal1 3710 326 3710 326 1 reg_six6
rlabel metal1 3710 318 3710 318 1 reg_six7
rlabel metal1 8013 2445 8013 2445 7 Y0
rlabel metal1 8012 2437 8012 2437 7 Y1
rlabel metal1 8012 2429 8012 2429 7 Y2
rlabel metal1 8011 2421 8011 2421 7 Y3
rlabel metal1 8012 2413 8012 2413 7 Y4
rlabel metal1 8012 2405 8012 2405 7 Y5
rlabel metal1 8012 2397 8012 2397 7 Y6
rlabel metal1 8013 2389 8013 2389 7 Y7
rlabel metal1 8012 2453 8012 2453 7 Overflow
rlabel metal1 8008 605 8008 605 1 Equal
rlabel metal2 3855 -10 3855 -10 1 RorL
rlabel metal3 96 3159 96 3159 1 VDD
rlabel metal3 163 -200 163 -200 1 VSS
rlabel m2contact 181 2610 181 2610 1 VDD
<< end >>
