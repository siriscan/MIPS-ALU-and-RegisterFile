magic
tech scmos
timestamp 1746219663
<< nwell >>
rect -8 39 97 92
<< ntransistor >>
rect 8 8 10 12
rect 18 8 20 12
rect 28 8 30 12
rect 38 8 40 12
rect 48 8 50 12
rect 58 8 60 12
rect 68 8 70 12
rect 78 8 80 12
<< ptransistor >>
rect 8 48 10 80
rect 18 48 20 80
rect 28 48 30 80
rect 38 48 40 80
rect 48 48 50 80
rect 58 48 60 80
rect 68 48 70 80
rect 78 48 80 80
<< ndiffusion >>
rect 6 8 8 12
rect 10 8 12 12
rect 16 8 18 12
rect 20 8 22 12
rect 26 8 28 12
rect 30 8 32 12
rect 36 8 38 12
rect 40 8 42 12
rect 46 8 48 12
rect 50 8 52 12
rect 56 8 58 12
rect 60 8 62 12
rect 66 8 68 12
rect 70 8 72 12
rect 76 8 78 12
rect 80 8 82 12
<< pdiffusion >>
rect 6 48 8 80
rect 10 48 18 80
rect 20 48 28 80
rect 30 48 38 80
rect 40 48 48 80
rect 50 48 58 80
rect 60 48 68 80
rect 70 48 78 80
rect 80 48 82 80
<< ndcontact >>
rect 2 8 6 12
rect 12 8 16 12
rect 22 8 26 12
rect 32 8 36 12
rect 42 8 46 12
rect 52 8 56 12
rect 62 8 66 12
rect 72 8 76 12
rect 82 8 86 12
<< pdcontact >>
rect 2 48 6 80
rect 82 48 86 80
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 84 6 88
<< polysilicon >>
rect 8 80 10 82
rect 18 80 20 82
rect 28 80 30 82
rect 38 80 40 82
rect 48 80 50 82
rect 58 80 60 82
rect 68 80 70 82
rect 78 80 80 82
rect 8 36 10 48
rect 18 36 20 48
rect 28 36 30 48
rect 38 36 40 48
rect 48 36 50 48
rect 58 36 60 48
rect 68 36 70 48
rect 78 36 80 48
rect 7 32 10 36
rect 17 32 20 36
rect 27 32 30 36
rect 37 32 40 36
rect 47 32 50 36
rect 57 32 60 36
rect 67 32 70 36
rect 77 32 80 36
rect 8 12 10 32
rect 18 12 20 32
rect 28 12 30 32
rect 38 12 40 32
rect 48 12 50 32
rect 58 12 60 32
rect 68 12 70 32
rect 78 12 80 32
rect 8 6 10 8
rect 18 6 20 8
rect 28 6 30 8
rect 38 6 40 8
rect 48 6 50 8
rect 58 6 60 8
rect 68 6 70 8
rect 78 6 80 8
<< polycontact >>
rect 3 32 7 36
rect 13 32 17 36
rect 23 32 27 36
rect 33 32 37 36
rect 43 32 47 36
rect 53 32 57 36
rect 63 32 67 36
rect 73 32 77 36
<< metal1 >>
rect 0 84 2 88
rect 6 84 88 88
rect 2 80 6 84
rect 82 24 86 48
rect 12 20 86 24
rect 12 12 16 20
rect 32 12 36 20
rect 52 12 56 20
rect 72 12 76 20
rect 2 4 6 8
rect 22 4 26 8
rect 42 4 46 8
rect 62 4 66 8
rect 82 4 86 8
rect 0 0 2 4
rect 6 0 88 4
<< labels >>
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel nsubstratencontact 4 86 4 86 1 VDD
rlabel polycontact 5 34 5 34 1 A
rlabel polycontact 15 34 15 34 1 B
rlabel polycontact 25 34 25 34 1 C
rlabel polycontact 35 34 35 34 1 D
rlabel polycontact 45 34 45 34 1 E
rlabel polycontact 55 34 55 34 1 F
rlabel polycontact 65 34 65 34 1 G
rlabel polycontact 75 34 75 34 1 H
rlabel metal1 84 32 84 32 1 Y
<< end >>
