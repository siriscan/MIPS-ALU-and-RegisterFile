magic
tech scmos
timestamp 1746070328
<< metal1 >>
rect -75 167 644 171
rect -67 159 833 163
rect -59 151 1023 155
rect -51 143 1214 147
rect -43 135 1402 139
rect -35 127 1591 131
rect -27 119 1781 123
rect -19 111 1972 115
rect 516 100 526 104
rect 516 16 526 20
rect -91 -8 54 -4
rect -91 -17 118 -13
rect -91 -25 182 -21
rect -91 -33 246 -29
rect -91 -41 310 -37
rect -91 -49 374 -45
rect -91 -57 438 -53
rect -91 -65 502 -61
rect 50 -78 543 -74
rect 114 -86 732 -82
rect 178 -94 922 -90
rect 242 -102 1113 -98
rect 306 -110 1301 -106
rect 370 -118 1490 -114
rect 434 -126 1680 -122
rect 498 -134 1871 -130
rect -19 -150 477 -146
rect -27 -158 413 -154
rect -35 -166 349 -162
rect -43 -174 285 -170
rect -51 -182 221 -178
rect -59 -190 157 -186
rect -67 -198 93 -194
rect -75 -206 29 -202
<< m2contact >>
rect -79 167 -75 171
rect 644 167 648 171
rect -71 159 -67 163
rect 833 159 837 163
rect -63 151 -59 155
rect 1023 151 1027 155
rect -55 143 -51 147
rect 1214 143 1218 147
rect -47 135 -43 139
rect 1402 135 1406 139
rect -39 127 -35 131
rect 1591 127 1595 131
rect -31 119 -27 123
rect 1781 119 1785 123
rect -23 111 -19 115
rect 1972 111 1976 115
rect 54 41 58 45
rect 118 40 122 44
rect 182 40 186 44
rect 246 39 250 43
rect 310 39 314 43
rect 374 41 378 45
rect 438 40 442 44
rect 502 40 506 44
rect 29 35 33 39
rect 93 31 97 35
rect 157 31 161 35
rect 221 31 225 35
rect 285 31 289 35
rect 349 31 353 35
rect 413 31 417 35
rect 477 31 481 35
rect 46 0 50 4
rect 110 0 114 4
rect 174 0 178 4
rect 238 0 242 4
rect 302 0 306 4
rect 366 0 370 4
rect 430 0 434 4
rect 494 0 498 4
rect 54 -8 58 -4
rect 118 -17 122 -13
rect 182 -25 186 -21
rect 246 -33 250 -29
rect 310 -41 314 -37
rect 374 -49 378 -45
rect 438 -57 442 -53
rect 502 -65 506 -61
rect 46 -78 50 -74
rect 543 -78 547 -74
rect 110 -86 114 -82
rect 732 -86 736 -82
rect 174 -94 178 -90
rect 922 -94 926 -90
rect 238 -102 242 -98
rect 1113 -102 1117 -98
rect 302 -110 306 -106
rect 1301 -110 1305 -106
rect 366 -118 370 -114
rect 1490 -118 1494 -114
rect 430 -126 434 -122
rect 1680 -126 1684 -122
rect 494 -134 498 -130
rect 1871 -134 1875 -130
rect -23 -150 -19 -146
rect 477 -150 481 -146
rect -31 -158 -27 -154
rect 413 -158 417 -154
rect -39 -166 -35 -162
rect 349 -166 353 -162
rect -47 -174 -43 -170
rect 285 -174 289 -170
rect -55 -182 -51 -178
rect 221 -182 225 -178
rect -63 -190 -59 -186
rect 157 -190 161 -186
rect -71 -198 -67 -194
rect 93 -198 97 -194
rect -79 -206 -75 -202
rect 29 -206 33 -202
<< metal2 >>
rect -79 -202 -75 167
rect -71 -194 -67 159
rect -63 -186 -59 151
rect -55 -178 -51 143
rect -47 -170 -43 135
rect -39 -162 -35 127
rect -31 -154 -27 119
rect -23 -146 -19 111
rect 6 -218 10 12
rect 29 -202 33 35
rect 46 -74 50 0
rect 54 -4 58 41
rect 93 -194 97 31
rect 110 -82 114 0
rect 118 -13 122 40
rect 157 -186 161 31
rect 174 -90 178 0
rect 182 -21 186 40
rect 221 -178 225 31
rect 238 -98 242 0
rect 246 -29 250 39
rect 285 -170 289 31
rect 302 -106 306 0
rect 310 -37 314 39
rect 349 -162 353 31
rect 366 -114 370 0
rect 374 -45 378 41
rect 413 -154 417 31
rect 430 -122 434 0
rect 438 -53 442 40
rect 477 -146 481 31
rect 494 -130 498 0
rect 502 -61 506 40
rect 543 -74 547 -32
rect 552 -218 556 12
rect 644 -218 648 167
rect 732 -82 736 -32
rect 833 -218 837 159
rect 922 -90 926 -32
rect 1023 -218 1027 151
rect 1113 -98 1117 -32
rect 1214 -218 1218 143
rect 1301 -106 1305 -31
rect 1402 -218 1406 135
rect 1490 -114 1494 -31
rect 1591 -218 1595 127
rect 1680 -122 1684 -32
rect 1781 -218 1785 119
rect 1871 -130 1875 -31
rect 1972 -218 1976 111
use reg8  reg8_0
timestamp 1745261002
transform 1 0 520 0 1 -16
box 0 -16 1512 124
use 8bitMUX2to1  8bitMUX2to1_0
timestamp 1746042099
transform 1 0 0 0 1 0
box 0 0 520 107
<< labels >>
rlabel metal1 518 113 518 113 1 A7
rlabel metal1 518 121 518 121 1 A6
rlabel metal1 518 129 518 129 1 A5
rlabel metal1 518 137 518 137 1 A4
rlabel metal1 518 145 518 145 1 A3
rlabel metal1 518 153 518 153 1 A2
rlabel metal1 518 161 518 161 1 A1
rlabel metal1 518 169 518 169 1 A0
rlabel metal1 521 18 521 18 1 VSS
rlabel metal1 520 102 521 102 1 VDD
rlabel metal1 2 -6 2 -6 1 D0
rlabel metal1 2 -15 2 -15 1 D1
rlabel metal1 2 -23 2 -23 1 D2
rlabel metal1 2 -31 2 -31 1 D3
rlabel metal1 2 -39 2 -39 1 D4
rlabel metal1 2 -47 2 -47 1 D5
rlabel metal1 2 -55 2 -55 1 D6
rlabel metal1 2 -63 2 -63 1 D7
rlabel metal2 8 -131 8 -131 1 EN
rlabel metal1 -89 -6 -89 -6 1 D0
rlabel metal1 -89 -15 -89 -15 1 D1
rlabel metal1 -89 -23 -89 -23 1 D2
rlabel metal1 -89 -31 -89 -31 1 D3
rlabel metal1 -89 -39 -89 -39 1 D4
rlabel metal1 -89 -47 -89 -47 1 D5
rlabel metal1 -89 -55 -89 -55 1 D6
rlabel metal1 -89 -63 -89 -63 1 D7
rlabel metal2 8 -216 8 -216 1 EN
rlabel metal2 554 -216 554 -216 1 CLK
rlabel metal2 1974 -216 1974 -216 1 Q7
rlabel metal2 1783 -216 1783 -216 1 Q6
rlabel metal2 1593 -216 1593 -216 1 Q5
rlabel metal2 1404 -216 1404 -216 1 Q4
rlabel metal2 1216 -216 1216 -216 1 Q3
rlabel metal2 1025 -216 1025 -216 1 Q2
rlabel metal2 835 -216 835 -216 1 Q1
rlabel metal2 646 -216 646 -216 1 Q0
<< end >>
